`timescale 1ns / 1ps
/*
	Input:
		时钟、复位
		din1, din2, din3, ...: 并行窗口数据
		df1_1, df1_2, df1_3, ...: 高斯滤波器参数，固定值
	Output:
		dout: 卷积结果输出
		out_en: 输出数据有效
	Description：
		功能上，2D卷积，将11x11窗口中的数据与卷积模块作乘积和操作；
		结构上，采用了11个一维卷积子模块，输入有11个88位的数据，分别表示窗口的11行，
		88位数据表示窗口一列11个8bit的数据，输入还有11个48位宽的模板参数，用于卷积。
		输出为18位宽的dout，为卷积结果。
	Note:
		由于高斯卷积的对称性，2D高斯卷积拆分成两个1D卷积，首先合并同类项，再去做乘法，减少DSP的使用数量。
		采用并行流水线结构，提高数据吞吐量
		在卷积运算过程中，需要对窗口数据做乘加操作，因此使用了Fuxi提供的内置DSP IP。
*/

module CONV(clk, rst, din1, din2, din3, din4, din5, din6, din7, din8, din9, din10, din11, 
				  df1_1, df1_2, df1_3, df1_4, df1_5, df1_6, df1_7, df1_8, df1_9, df1_10, df1_11,
				  dout,out_en);
    input clk;
    input rst;
    input [87:0] din1;
    input [87:0] din2;
    input [87:0] din3;
    input [87:0] din4;
    input [87:0] din5;
    input [87:0] din6;
    input [87:0] din7;
    input [87:0] din8;
    input [87:0] din9;
    input [87:0] din10;
    input [87:0] din11;
	 
	input [47:0] df1_1;
	input [47:0] df1_2;
	input [47:0] df1_3;
	input [47:0] df1_4;
	input [47:0] df1_5;
	input [47:0] df1_6;
	input [47:0] df1_7;
	input [47:0] df1_8;
	input [47:0] df1_9;
	input [47:0] df1_10;
	input [47:0] df1_11;
	 
    output [17:0] dout;
    output out_en;
	 
	 //**********************输出赋值 ******************************//
	reg [23:0] dout1;
	wire [17:0] dout;  reg [4:0] cnt_out_en; reg out_en;
	assign dout=dout1[17:0];
	
	always @(posedge clk or negedge rst)
	begin
	if(!rst)
	begin
		out_en<=0;
		cnt_out_en<=0;
	end
	else
	begin
		if(cnt_out_en>=10)
			out_en<=1;
		else
		begin
			cnt_out_en<=cnt_out_en+1;
			out_en<=0;
		end
	end
	end
	
	//*****************  图像数据  *******************************//	
	wire [7:0] d1[10:0];wire [7:0] d2[10:0];wire [7:0] d3[10:0];wire [7:0] d4[10:0];wire [7:0] d5[10:0];
	wire [7:0] d6[10:0];wire [7:0] d7[10:0];wire [7:0] d8[10:0];wire [7:0] d9[10:0];wire [7:0] d10[10:0];
	wire [7:0] d11[10:0];

	//****************   DoG  参数   ****************************// 
	wire [7:0] k1_1[5:0];wire [7:0] k1_2[5:0];wire [7:0] k1_3[5:0];wire [7:0] k1_4[5:0];wire [7:0] k1_5[5:0];
	wire [7:0] k1_6[5:0];wire [7:0] k1_7[5:0];wire [7:0] k1_8[5:0];wire [7:0] k1_9[5:0];wire [7:0] k1_10[5:0];
	wire [7:0] k1_11[5:0];

	// ***************** 图像数据赋值************************//
	assign {d1[10],d1[9],d1[8],d1[7],d1[6],d1[5],d1[4],d1[3],d1[2],d1[1],d1[0]}=din1;
	assign {d2[10],d2[9],d2[8],d2[7],d2[6],d2[5],d2[4],d2[3],d2[2],d2[1],d2[0]}=din2;
	assign {d3[10],d3[9],d3[8],d3[7],d3[6],d3[5],d3[4],d3[3],d3[2],d3[1],d3[0]}=din3;
	assign {d4[10],d4[9],d4[8],d4[7],d4[6],d4[5],d4[4],d4[3],d4[2],d4[1],d4[0]}=din4;
	assign {d5[10],d5[9],d5[8],d5[7],d5[6],d5[5],d5[4],d5[3],d5[2],d5[1],d5[0]}=din5;
	assign {d6[10],d6[9],d6[8],d6[7],d6[6],d6[5],d6[4],d6[3],d6[2],d6[1],d6[0]}=din6;
	assign {d7[10],d7[9],d7[8],d7[7],d7[6],d7[5],d7[4],d7[3],d7[2],d7[1],d7[0]}=din7;
	assign {d8[10],d8[9],d8[8],d8[7],d8[6],d8[5],d8[4],d8[3],d8[2],d8[1],d8[0]}=din8;
	assign {d9[10],d9[9],d9[8],d9[7],d9[6],d9[5],d9[4],d9[3],d9[2],d9[1],d9[0]}=din9;
	assign {d10[10],d10[9],d10[8],d10[7],d10[6],d10[5],d10[4],d10[3],d10[2],d10[1],d10[0]}=din10;
	assign {d11[10],d11[9],d11[8],d11[7],d11[6],d11[5],d11[4],d11[3],d11[2],d11[1],d11[0]}=din11;

 //********************* DoG 参数赋值 **************************//
	assign {k1_1[5],k1_1[4],k1_1[3],k1_1[2],k1_1[1],k1_1[0]}=df1_1;
	assign {k1_2[5],k1_2[4],k1_2[3],k1_2[2],k1_2[1],k1_2[0]}=df1_2;
	assign {k1_3[5],k1_3[4],k1_3[3],k1_3[2],k1_3[1],k1_3[0]}=df1_3;
	assign {k1_4[5],k1_4[4],k1_4[3],k1_4[2],k1_4[1],k1_4[0]}=df1_4;
	assign {k1_5[5],k1_5[4],k1_5[3],k1_5[2],k1_5[1],k1_5[0]}=df1_5;
	assign {k1_6[5],k1_6[4],k1_6[3],k1_6[2],k1_6[1],k1_6[0]}=df1_6;
	assign {k1_7[5],k1_7[4],k1_7[3],k1_7[2],k1_7[1],k1_7[0]}=df1_7;
	assign {k1_8[5],k1_8[4],k1_8[3],k1_8[2],k1_8[1],k1_8[0]}=df1_8;
	assign {k1_9[5],k1_9[4],k1_9[3],k1_9[2],k1_9[1],k1_9[0]}=df1_9;
	assign {k1_10[5],k1_10[4],k1_10[3],k1_10[2],k1_10[1],k1_10[0]}=df1_10;
	assign {k1_11[5],k1_11[4],k1_11[3],k1_11[2],k1_11[1],k1_11[0]}=df1_11;

	
	//**********************************  卷积运算  ***********************//
	wire [20:0] r1_1[4:0];
	reg [21:0] r1_2[2:0];
	reg [22:0] r1_3[1:0];

	reg [8:0] ra1_1[5:0];
	reg [8:0] ra1_2[5:0];
	reg [8:0] ra1_3[5:0];
	reg [8:0] ra1_4[5:0];
	reg [8:0] ra1_5[5:0];
	reg [8:0] ra1_6[5:0];
	reg [8:0] ra1_7[5:0];
	reg [8:0] ra1_8[5:0];
	reg [8:0] ra1_9[5:0];
	reg [8:0] ra1_10[5:0];
	reg [8:0] ra1_11[5:0];
	
	reg [9:0] ra2_1[5:0];
	reg [9:0] ra2_2[5:0];
	reg [9:0] ra2_3[5:0];
	reg [9:0] ra2_4[5:0];
	reg [9:0] ra2_5[5:0];
	reg [9:0] ra2_6[5:0];
	 
	//*******************************卷积————加法运算 ************************//
	always @(posedge clk,negedge rst)
	begin
		if(!rst)
		begin
			dout1 <= 'd0;
		end
		else
		begin
	//*************		对称加法	************* //
			ra1_1[0]<=d1[0]+d1[10];ra1_1[2]<=d1[2]+d1[8];ra1_1[4]<=d1[4]+d1[6];
			ra1_1[1]<=d1[1]+d1[9]; ra1_1[3]<=d1[3]+d1[7];ra1_1[5]<=d1[5];
			
			ra1_2[0]<=d2[0]+d2[10];ra1_2[2]<=d2[2]+d2[8];ra1_2[4]<=d2[4]+d2[6];
			ra1_2[1]<=d2[1]+d2[9]; ra1_2[3]<=d2[3]+d2[7];ra1_2[5]<=d2[5];
			
			ra1_3[0]<=d3[0]+d3[10];ra1_3[2]<=d3[2]+d3[8];ra1_3[4]<=d3[4]+d3[6];
			ra1_3[1]<=d3[1]+d3[9]; ra1_3[3]<=d3[3]+d3[7];ra1_3[5]<=d3[5];
			
			ra1_4[0]<=d4[0]+d4[10];ra1_4[2]<=d4[2]+d4[8];ra1_4[4]<=d4[4]+d4[6];
			ra1_4[1]<=d4[1]+d4[9]; ra1_4[3]<=d4[3]+d4[7];ra1_4[5]<=d4[5];
			
			ra1_5[0]<=d5[0]+d5[10];ra1_5[2]<=d5[2]+d5[8];ra1_5[4]<=d5[4]+d5[6];
			ra1_5[1]<=d5[1]+d5[9]; ra1_5[3]<=d5[3]+d5[7];ra1_5[5]<=d5[5];
			
			ra1_6[0]<=d6[0]+d6[10];ra1_6[2]<=d6[2]+d6[8];ra1_6[4]<=d6[4]+d6[6];
			ra1_6[1]<=d6[1]+d6[9]; ra1_6[3]<=d6[3]+d6[7];ra1_6[5]<=d6[5];
			
			ra1_7[0]<=d7[0]+d7[10];ra1_7[2]<=d7[2]+d7[8];ra1_7[4]<=d7[4]+d7[6];
			ra1_7[1]<=d7[1]+d7[9]; ra1_7[3]<=d7[3]+d7[7];ra1_7[5]<=d7[5];
			
			ra1_8[0]<=d8[0]+d8[10];ra1_8[2]<=d8[2]+d8[8];ra1_8[4]<=d8[4]+d8[6];
			ra1_8[1]<=d8[1]+d8[9]; ra1_8[3]<=d8[3]+d8[7];ra1_8[5]<=d8[5];
			
			ra1_9[0]<=d9[0]+d9[10];ra1_9[2]<=d9[2]+d9[8];ra1_9[4]<=d9[4]+d9[6];
			ra1_9[1]<=d9[1]+d9[9]; ra1_9[3]<=d9[3]+d9[7];ra1_9[5]<=d9[5];
			
			ra1_10[0]<=d10[0]+d10[10];ra1_10[2]<=d10[2]+d10[8];ra1_10[4]<=d10[4]+d10[6];
			ra1_10[1]<=d10[1]+d10[9]; ra1_10[3]<=d10[3]+d10[7];ra1_10[5]<=d10[5];
			
			ra1_11[0]<=d11[0]+d11[10];ra1_11[2]<=d11[2]+d11[8];ra1_11[4]<=d11[4]+d11[6];
			ra1_11[1]<=d11[1]+d11[9]; ra1_11[3]<=d11[3]+d11[7];ra1_11[5]<=d11[5];
			
			ra2_1[0]<=ra1_1[0]+ra1_11[0];ra2_1[2]<=ra1_1[2]+ra1_11[2];ra2_1[4]<=ra1_1[4]+ra1_11[4];
			ra2_1[1]<=ra1_1[1]+ra1_11[1];ra2_1[3]<=ra1_1[3]+ra1_11[3];ra2_1[5]<=ra1_1[5]+ra1_11[5];
			
			ra2_2[0]<=ra1_2[0]+ra1_10[0];ra2_2[2]<=ra1_2[2]+ra1_10[2];ra2_2[4]<=ra1_2[4]+ra1_10[4];
			ra2_2[1]<=ra1_2[1]+ra1_10[1];ra2_2[3]<=ra1_2[3]+ra1_10[3];ra2_2[5]<=ra1_2[5]+ra1_10[5];
			
			ra2_3[0]<=ra1_3[0]+ra1_9[0];ra2_3[2]<=ra1_3[2]+ra1_9[2];ra2_3[4]<=ra1_3[4]+ra1_9[4];
			ra2_3[1]<=ra1_3[1]+ra1_9[1];ra2_3[3]<=ra1_3[3]+ra1_9[3];ra2_3[5]<=ra1_3[5]+ra1_9[5];			
			
			ra2_4[0]<=ra1_4[0]+ra1_8[0];ra2_4[2]<=ra1_4[2]+ra1_8[2];ra2_4[4]<=ra1_4[4]+ra1_8[4];
			ra2_4[1]<=ra1_4[1]+ra1_8[1];ra2_4[3]<=ra1_4[3]+ra1_8[3];ra2_4[5]<=ra1_4[5]+ra1_8[5];

			ra2_5[0]<=ra1_5[0]+ra1_7[0];ra2_5[2]<=ra1_5[2]+ra1_7[2];ra2_5[4]<=ra1_5[4]+ra1_7[4];
			ra2_5[1]<=ra1_5[1]+ra1_7[1];ra2_5[3]<=ra1_5[3]+ra1_7[3];ra2_5[5]<=ra1_5[5]+ra1_7[5];

			ra2_6[0]<=ra1_6[0];ra2_6[2]<=ra1_6[2];ra2_6[4]<=ra1_6[4];
			ra2_6[1]<=ra1_6[1];ra2_6[3]<=ra1_6[3];ra2_6[5]<=ra1_6[5];			
			
	//**************乘法结果做加法
			
			r1_2[0]<=r1_1[0]+r1_1[4];
			r1_2[1]<=r1_1[1]+r1_1[3];
			r1_2[2]<=r1_1[2];	
			r1_3[0]<=r1_2[0]+r1_2[1];
			r1_3[1]<=r1_2[2];
	
			dout1<=r1_3[0]+r1_3[1];
		end
	end
	 
	 
	 //************************ 卷积————乘加运算*********************//
	cov cov1_1(
		.clk(clk), .rst(rst), 
		
		.din1(ra2_1[0]), .din2(ra2_1[1]), .din3(ra2_1[2]), .din4(ra2_1[3]), 
		.din5(ra2_1[4]), .din6(ra2_1[5]),.din7(ra2_2[0]), .din8(ra2_2[1]),
	
		.k1(k1_1[5]), .k2(k1_1[4]), .k3(k1_1[3]),.k4(k1_1[2]),.k5(k1_1[1]), 
		.k6(k1_1[0]), .k7(k1_2[5]), .k8(k1_2[4]),
		.dout(r1_1[0])
	);
	
	
				  
	cov cov1_2(
		.clk(clk), .rst(rst),  
		
		.din1(ra2_2[2]), .din2(ra2_2[3]), .din3(ra2_2[4]), .din4(ra2_2[5]), 
		.din5(ra2_3[0]), .din6(ra2_3[1]), .din7(ra2_3[2]), .din8(ra2_3[3]),
		
		.k1(k1_2[3]), .k2(k1_2[2]), .k3(k1_2[1]),.k4(k1_2[0]),.k5(k1_3[5]), 
		.k6(k1_3[4]), .k7(k1_3[3]), .k8(k1_3[2]),
		.dout(r1_1[1])
	);
				  
				  
	cov cov1_3(	  
		.clk(clk), .rst(rst),  
		
		.din1(ra2_3[4]), .din2(ra2_3[5]), .din3(ra2_4[0]), .din4(ra2_4[1]),
		.din5(ra2_4[2]), .din6(ra2_4[3]), .din7(ra2_4[4]), .din8(ra2_4[5]),
				  
		.k1(k1_3[1]), .k2(k1_3[0]), .k3(k1_4[5]),.k4(k1_4[4]),.k5(k1_4[3]),
		.k6(k1_4[2]), .k7(k1_4[1]), .k8(k1_4[0]),
				  
		.dout(r1_1[2])
	);
				  
				  
				  
	cov cov1_4(
		.clk(clk), .rst(rst), 
	
		.din1(ra2_5[0]), .din2(ra2_5[1]), .din3(ra2_5[2]), .din4(ra2_5[3]),
		.din5(ra2_5[4]), .din6(ra2_5[5]),.din7(ra2_6[0]), .din8(ra2_6[1]),
				  
		.k1(k1_5[5]), .k2(k1_5[4]), .k3(k1_5[3]),.k4(k1_5[2]),.k5(k1_5[1]),
		.k6(k1_5[0]), .k7(k1_6[5]), .k8(k1_6[4]),
				  
		.dout(r1_1[3])
	);
				  
				  		  
	cov cov1_5(
		.clk(clk), .rst(rst), 
		
		.din1(ra2_6[2]), .din2(ra2_6[3]), .din3(ra2_6[4]), .din4(ra2_6[5]),
		.din5(0), .din6(0),.din7(0), .din8(0),
		
		.k1(k1_6[3]), .k2(k1_6[2]), .k3(k1_6[1]),.k4(k1_6[0]),.k5(0),
		.k6(0), .k7(0), .k8(0),

		.dout(r1_1[4])
	);
				  

	
endmodule
