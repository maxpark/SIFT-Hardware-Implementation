`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:34:16 06/13/2022 
// Design Name: 
// Module Name:    dir34_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module dir34_1
(
    input   [7:0]       a,  // Addr.
	output  reg [4:0]	spo // Data.
);
	
	always @(*) begin
		case (a)
			000: spo = 5'h16;
            001: spo = 5'h16;
            002: spo = 5'h16;
            003: spo = 5'h17;
            004: spo = 5'h17;
            005: spo = 5'h17;
            006: spo = 5'h18;
            007: spo = 5'h18;
            008: spo = 5'h18;
            009: spo = 5'h19;
            010: spo = 5'h19;
            011: spo = 5'h1a;
            012: spo = 5'h1a;
            013: spo = 5'h1a;
            014: spo = 5'h1b;
            015: spo = 5'h1b;
            016: spo = 5'h17;
            017: spo = 5'h17;
            018: spo = 5'h17;
            019: spo = 5'h18;
            020: spo = 5'h18;
            021: spo = 5'h18;
            022: spo = 5'h19;
            023: spo = 5'h19;
            024: spo = 5'h19;
            025: spo = 5'h1a;
            026: spo = 5'h1a;
            027: spo = 5'h1a;
            028: spo = 5'h1b;
            029: spo = 5'h1b;
            030: spo = 5'h1b;
            031: spo = 5'h1c;
            032: spo = 5'h18;
            033: spo = 5'h18;
            034: spo = 5'h18;
            035: spo = 5'h19;
            036: spo = 5'h19;
            037: spo = 5'h19;
            038: spo = 5'h1a;
            039: spo = 5'h1a;
            040: spo = 5'h1a;
            041: spo = 5'h1b;
            042: spo = 5'h1b;
            043: spo = 5'h1b;
            044: spo = 5'h1c;
            045: spo = 5'h1c;
            046: spo = 5'h1c;
            047: spo = 5'h1d;
            048: spo = 5'h19;
            049: spo = 5'h19;
            050: spo = 5'h19;
            051: spo = 5'h1a;
            052: spo = 5'h1a;
            053: spo = 5'h1a;
            054: spo = 5'h1b;
            055: spo = 5'h1b;
            056: spo = 5'h1b;
            057: spo = 5'h1c;
            058: spo = 5'h1c;
            059: spo = 5'h1c;
            060: spo = 5'h1d;
            061: spo = 5'h1d;
            062: spo = 5'h1d;
            063: spo = 5'h1e;
            064: spo = 5'h1a;
            065: spo = 5'h1a;
            066: spo = 5'h1a;
            067: spo = 5'h1b;
            068: spo = 5'h1b;
            069: spo = 5'h1b;
            070: spo = 5'h1c;
            071: spo = 5'h1c;
            072: spo = 5'h1c;
            073: spo = 5'h1d;
            074: spo = 5'h1d;
            075: spo = 5'h1d;
            076: spo = 5'h1e;
            077: spo = 5'h1e;
            078: spo = 5'h1e;
            079: spo = 5'h1f;
            080: spo = 5'h1a;
            081: spo = 5'h1b;
            082: spo = 5'h1b;
            083: spo = 5'h1b;
            084: spo = 5'h1c;
            085: spo = 5'h1c;
            086: spo = 5'h1c;
            087: spo = 5'h1d;
            088: spo = 5'h1d;
            089: spo = 5'h1e;
            090: spo = 5'h1e;
            091: spo = 5'h1e;
            092: spo = 5'h1f;
            093: spo = 5'h1f;
            094: spo = 5'h1f;
            095: spo = 5'h0;
            096: spo = 5'h1b;
            097: spo = 5'h1c;
            098: spo = 5'h1c;
            099: spo = 5'h1c;
            100: spo = 5'h1d;
            101: spo = 5'h1d;
            102: spo = 5'h1d;
            103: spo = 5'h1e;
            104: spo = 5'h1e;
            105: spo = 5'h1e;
            106: spo = 5'h1f;
            107: spo = 5'h1f;
            108: spo = 5'h1f;
            109: spo = 5'h0;
            110: spo = 5'h0;
            111: spo = 5'h1;
            112: spo = 5'h1c;
            113: spo = 5'h1d;
            114: spo = 5'h1d;
            115: spo = 5'h1d;
            116: spo = 5'h1e;
            117: spo = 5'h1e;
            118: spo = 5'h1e;
            119: spo = 5'h1f;
            120: spo = 5'h1f;
            121: spo = 5'h1f;
            122: spo = 5'h0;
            123: spo = 5'h0;
            124: spo = 5'h0;
            125: spo = 5'h1;
            126: spo = 5'h1;
            127: spo = 5'h1;
            128: spo = 5'h1d;
            129: spo = 5'h1e;
            130: spo = 5'h1e;
            131: spo = 5'h1e;
            132: spo = 5'h1f;
            133: spo = 5'h1f;
            134: spo = 5'h1f;
            135: spo = 5'h0;
            136: spo = 5'h0;
            137: spo = 5'h0;
            138: spo = 5'h1;
            139: spo = 5'h1;
            140: spo = 5'h1;
            141: spo = 5'h2;
            142: spo = 5'h2;
            143: spo = 5'h2;
            144: spo = 5'h1e;
            145: spo = 5'h1f;
            146: spo = 5'h1f;
            147: spo = 5'h1f;
            148: spo = 5'h0;
            149: spo = 5'h0;
            150: spo = 5'h0;
            151: spo = 5'h1;
            152: spo = 5'h1;
            153: spo = 5'h1;
            154: spo = 5'h2;
            155: spo = 5'h2;
            156: spo = 5'h2;
            157: spo = 5'h3;
            158: spo = 5'h3;
            159: spo = 5'h3;
            160: spo = 5'h1f;
            161: spo = 5'h1f;
            162: spo = 5'h0;
            163: spo = 5'h0;
            164: spo = 5'h1;
            165: spo = 5'h1;
            166: spo = 5'h1;
            167: spo = 5'h2;
            168: spo = 5'h2;
            169: spo = 5'h2;
            170: spo = 5'h3;
            171: spo = 5'h3;
            172: spo = 5'h3;
            173: spo = 5'h4;
            174: spo = 5'h4;
            175: spo = 5'h4;
            176: spo = 5'h0;
            177: spo = 5'h0;
            178: spo = 5'h1;
            179: spo = 5'h1;
            180: spo = 5'h1;
            181: spo = 5'h2;
            182: spo = 5'h2;
            183: spo = 5'h2;
            184: spo = 5'h3;
            185: spo = 5'h3;
            186: spo = 5'h4;
            187: spo = 5'h4;
            188: spo = 5'h4;
            189: spo = 5'h5;
            190: spo = 5'h5;
            191: spo = 5'h5;
            192: spo = 5'h1;
            193: spo = 5'h1;
            194: spo = 5'h2;
            195: spo = 5'h2;
            196: spo = 5'h2;
            197: spo = 5'h3;
            198: spo = 5'h3;
            199: spo = 5'h3;
            200: spo = 5'h4;
            201: spo = 5'h4;
            202: spo = 5'h4;
            203: spo = 5'h5;
            204: spo = 5'h5;
            205: spo = 5'h5;
            206: spo = 5'h6;
            207: spo = 5'h6;
            208: spo = 5'h2;
            209: spo = 5'h2;
            210: spo = 5'h3;
            211: spo = 5'h3;
            212: spo = 5'h3;
            213: spo = 5'h4;
            214: spo = 5'h4;
            215: spo = 5'h4;
            216: spo = 5'h5;
            217: spo = 5'h5;
            218: spo = 5'h5;
            219: spo = 5'h6;
            220: spo = 5'h6;
            221: spo = 5'h6;
            222: spo = 5'h7;
            223: spo = 5'h7;
            224: spo = 5'h3;
            225: spo = 5'h3;
            226: spo = 5'h4;
            227: spo = 5'h4;
            228: spo = 5'h4;
            229: spo = 5'h5;
            230: spo = 5'h5;
            231: spo = 5'h5;
            232: spo = 5'h6;
            233: spo = 5'h6;
            234: spo = 5'h6;
            235: spo = 5'h7;
            236: spo = 5'h7;
            237: spo = 5'h7;
            238: spo = 5'h8;
            239: spo = 5'h8;
            240: spo = 5'h4;
            241: spo = 5'h4;
            242: spo = 5'h5;
            243: spo = 5'h5;
            244: spo = 5'h5;
            245: spo = 5'h6;
            246: spo = 5'h6;
            247: spo = 5'h6;
            248: spo = 5'h7;
            249: spo = 5'h7;
            250: spo = 5'h7;
            251: spo = 5'h8;
            252: spo = 5'h8;
            253: spo = 5'h8;
            254: spo = 5'h9;
            255: spo = 5'h9;
            default: spo = 5'h0;
		endcase
	end
endmodule