module fifo2ram_emb_v1 (clkr, clkw, cer, cew, rstnr, ar, aw, dw, qr);
input clkr;
input clkw;
input cer;
input cew;
input rstnr;
input [17:0] ar;
input [13:0] aw;
input [127:0] dw;
output [7:0] qr;

wire vcc_net;
wire gnd_net;
wire net_3;
wire net_33;
wire net_35;
wire net_36;
wire net_37;
wire addra_pipe_0_net;
wire net_41;
wire net_42;
wire net_43;
wire net_44;
wire net_45;
wire net_46;
wire net_48;
wire net_49;
wire net_50;
wire net_52;
wire net_53;
wire net_54;
wire addra_pipe_1_net;
wire net_56;
wire net_57;
wire net_58;
wire net_59;
wire net_60;
wire net_61;
wire net_63;
wire net_64;
wire net_65;
wire net_67;
wire net_68;
wire net_69;
wire net_70;
wire net_71;
wire net_72;
wire net_74;
wire net_75;
wire net_76;
wire net_78;
wire net_79;
wire net_80;
wire net_81;
wire net_82;
wire net_83;
wire addra_pipe_2_net;
wire net_85;
wire net_86;
wire net_87;
wire net_88;
wire net_89;
wire net_90;
wire net_92;
wire net_93;
wire net_94;
wire net_96;
wire net_97;
wire net_98;
wire net_99;
wire net_100;
wire net_101;
wire net_103;
wire net_104;
wire net_105;
wire net_107;
wire net_108;
wire net_109;
wire net_110;
wire net_111;
wire net_112;
wire net_113;
wire net_114;
wire net_115;
wire net_117;
wire net_118;
wire net_119;
wire net_121;
wire net_122;
wire net_123;
wire net_124;
wire net_125;
wire net_126;
wire net_128;
wire net_129;
wire net_130;
wire net_132;
wire net_133;
wire net_134;
wire net_135;
wire net_136;
wire net_137;
wire net_138;
wire net_139;
wire net_140;
wire addra_pipe_3_net;
wire net_143;
wire net_145;
wire net_146;
wire net_147;
wire net_149;
wire net_150;
wire net_151;
wire net_153;
wire net_154;
wire net_155;
wire net_156;
wire net_157;
wire net_158;
wire net_160;
wire net_161;
wire net_162;
wire net_164;
wire net_165;
wire net_166;
wire net_167;
wire net_168;
wire net_169;
wire net_170;
wire net_171;
wire net_172;
wire net_174;
wire net_175;
wire net_176;
wire net_178;
wire net_179;
wire net_180;
wire net_181;
wire net_182;
wire net_183;
wire net_185;
wire net_186;
wire net_187;
wire net_189;
wire net_190;
wire net_191;
wire net_192;
wire net_193;
wire net_194;
wire net_195;
wire net_196;
wire net_197;
wire net_198;
wire net_199;
wire net_200;
wire net_202;
wire net_203;
wire net_204;
wire net_206;
wire net_207;
wire net_208;
wire net_209;
wire net_210;
wire net_211;
wire net_213;
wire net_214;
wire net_215;
wire net_217;
wire net_218;
wire net_219;
wire net_220;
wire net_221;
wire net_222;
wire net_223;
wire net_224;
wire net_225;
wire net_227;
wire net_228;
wire net_229;
wire net_231;
wire net_232;
wire net_233;
wire net_234;
wire net_235;
wire net_236;
wire net_238;
wire net_239;
wire net_240;
wire net_242;
wire net_243;
wire net_244;
wire net_245;
wire net_246;
wire net_247;
wire net_248;
wire net_249;
wire net_250;
wire net_252;
wire net_253;
wire net_254;
wire net_255;
wire net_256;
wire net_258;
wire net_259;
wire net_260;
wire net_262;
wire net_263;
wire net_264;
wire net_265;
wire net_266;
wire net_267;
wire net_269;
wire net_270;
wire net_271;
wire net_273;
wire net_274;
wire net_275;
wire net_276;
wire net_277;
wire net_278;
wire net_279;
wire net_280;
wire net_281;
wire net_283;
wire net_284;
wire net_285;
wire net_287;
wire net_288;
wire net_289;
wire net_290;
wire net_291;
wire net_292;
wire net_294;
wire net_295;
wire net_296;
wire net_298;
wire net_299;
wire net_300;
wire net_301;
wire net_302;
wire net_303;
wire net_304;
wire net_305;
wire net_306;
wire net_307;
wire net_308;
wire net_309;
wire net_311;
wire net_312;
wire net_313;
wire net_315;
wire net_316;
wire net_317;
wire net_318;
wire net_319;
wire net_320;
wire net_322;
wire net_323;
wire net_324;
wire net_326;
wire net_327;
wire net_328;
wire net_329;
wire net_330;
wire net_331;
wire net_332;
wire net_333;
wire net_334;
wire net_336;
wire net_337;
wire net_338;
wire net_340;
wire net_341;
wire net_342;
wire net_343;
wire net_344;
wire net_345;
wire net_347;
wire net_348;
wire net_349;
wire net_351;
wire net_352;
wire net_353;
wire net_354;
wire net_355;
wire net_356;
wire net_357;
wire net_358;
wire net_359;
wire net_361;
wire net_362;
wire net_363;
wire net_364;
wire net_365;
wire net_367;
wire net_368;
wire net_369;
wire net_371;
wire net_372;
wire net_373;
wire net_374;
wire net_375;
wire net_376;
wire net_378;
wire net_379;
wire net_380;
wire net_382;
wire net_383;
wire net_384;
wire net_385;
wire net_386;
wire net_387;
wire net_388;
wire net_389;
wire net_390;
wire net_392;
wire net_393;
wire net_394;
wire net_396;
wire net_397;
wire net_398;
wire net_399;
wire net_400;
wire net_401;
wire net_403;
wire net_404;
wire net_405;
wire net_407;
wire net_408;
wire net_409;
wire net_410;
wire net_411;
wire net_412;
wire net_413;
wire net_414;
wire net_415;
wire net_416;
wire net_417;
wire net_418;
wire net_420;
wire net_421;
wire net_422;
wire net_424;
wire net_425;
wire net_426;
wire net_427;
wire net_428;
wire net_429;
wire net_431;
wire net_432;
wire net_433;
wire net_435;
wire net_436;
wire net_437;
wire net_438;
wire net_439;
wire net_440;
wire net_441;
wire net_442;
wire net_443;
wire net_445;
wire net_446;
wire net_447;
wire net_449;
wire net_450;
wire net_451;
wire net_452;
wire net_453;
wire net_454;
wire net_456;
wire net_457;
wire net_458;
wire net_460;
wire net_461;
wire net_462;
wire net_463;
wire net_464;
wire net_465;
wire net_466;
wire net_467;
wire net_468;
wire net_470;
wire net_471;
wire net_472;
wire net_473;
wire net_474;
wire net_476;
wire net_477;
wire net_478;
wire net_480;
wire net_481;
wire net_482;
wire net_483;
wire net_484;
wire net_485;
wire net_487;
wire net_488;
wire net_489;
wire net_491;
wire net_492;
wire net_493;
wire net_494;
wire net_495;
wire net_496;
wire net_497;
wire net_498;
wire net_499;
wire net_501;
wire net_502;
wire net_503;
wire net_505;
wire net_506;
wire net_507;
wire net_508;
wire net_509;
wire net_510;
wire net_512;
wire net_513;
wire net_514;
wire net_516;
wire net_517;
wire net_518;
wire net_519;
wire net_520;
wire net_521;
wire net_522;
wire net_523;
wire net_524;
wire net_525;
wire net_526;
wire net_527;
wire net_529;
wire net_530;
wire net_531;
wire net_533;
wire net_534;
wire net_535;
wire net_536;
wire net_537;
wire net_538;
wire net_540;
wire net_541;
wire net_542;
wire net_544;
wire net_545;
wire net_546;
wire net_547;
wire net_548;
wire net_549;
wire net_550;
wire net_551;
wire net_552;
wire net_554;
wire net_555;
wire net_556;
wire net_558;
wire net_559;
wire net_560;
wire net_561;
wire net_562;
wire net_563;
wire net_565;
wire net_566;
wire net_567;
wire net_569;
wire net_570;
wire net_571;
wire net_572;
wire net_573;
wire net_574;
wire net_575;
wire net_576;
wire net_577;
wire net_579;
wire net_580;
wire net_581;
wire net_582;
wire net_583;
wire net_585;
wire net_586;
wire net_587;
wire net_589;
wire net_590;
wire net_591;
wire net_592;
wire net_593;
wire net_594;
wire net_596;
wire net_597;
wire net_598;
wire net_600;
wire net_601;
wire net_602;
wire net_603;
wire net_604;
wire net_605;
wire net_606;
wire net_607;
wire net_608;
wire net_610;
wire net_611;
wire net_612;
wire net_614;
wire net_615;
wire net_616;
wire net_617;
wire net_618;
wire net_619;
wire net_621;
wire net_622;
wire net_623;
wire net_625;
wire net_626;
wire net_627;
wire net_628;
wire net_629;
wire net_630;
wire net_631;
wire net_632;
wire net_633;
wire net_634;
wire net_635;
wire net_636;
wire net_638;
wire net_639;
wire net_640;
wire net_642;
wire net_643;
wire net_644;
wire net_645;
wire net_646;
wire net_647;
wire net_649;
wire net_650;
wire net_651;
wire net_653;
wire net_654;
wire net_655;
wire net_656;
wire net_657;
wire net_658;
wire net_659;
wire net_660;
wire net_661;
wire net_663;
wire net_664;
wire net_665;
wire net_667;
wire net_668;
wire net_669;
wire net_670;
wire net_671;
wire net_672;
wire net_674;
wire net_675;
wire net_676;
wire net_678;
wire net_679;
wire net_680;
wire net_681;
wire net_682;
wire net_683;
wire net_684;
wire net_685;
wire net_686;
wire net_688;
wire net_689;
wire net_690;
wire net_691;
wire net_692;
wire net_694;
wire net_695;
wire net_696;
wire net_698;
wire net_699;
wire net_700;
wire net_701;
wire net_702;
wire net_703;
wire net_705;
wire net_706;
wire net_707;
wire net_709;
wire net_710;
wire net_711;
wire net_712;
wire net_713;
wire net_714;
wire net_715;
wire net_716;
wire net_717;
wire net_719;
wire net_720;
wire net_721;
wire net_723;
wire net_724;
wire net_725;
wire net_726;
wire net_727;
wire net_728;
wire net_730;
wire net_731;
wire net_732;
wire net_734;
wire net_735;
wire net_736;
wire net_737;
wire net_738;
wire net_739;
wire net_740;
wire net_741;
wire net_742;
wire net_743;
wire net_744;
wire net_745;
wire net_747;
wire net_748;
wire net_749;
wire net_751;
wire net_752;
wire net_753;
wire net_754;
wire net_755;
wire net_756;
wire net_758;
wire net_759;
wire net_760;
wire net_762;
wire net_763;
wire net_764;
wire net_765;
wire net_766;
wire net_767;
wire net_768;
wire net_769;
wire net_770;
wire net_772;
wire net_773;
wire net_774;
wire net_776;
wire net_777;
wire net_778;
wire net_779;
wire net_780;
wire net_781;
wire net_783;
wire net_784;
wire net_785;
wire net_787;
wire net_788;
wire net_789;
wire net_790;
wire net_791;
wire net_792;
wire net_793;
wire net_794;
wire net_795;
wire net_797;
wire net_798;
wire net_799;
wire net_800;
wire net_801;
wire net_803;
wire net_804;
wire net_805;
wire net_807;
wire net_808;
wire net_809;
wire net_810;
wire net_811;
wire net_812;
wire net_814;
wire net_815;
wire net_816;
wire net_818;
wire net_819;
wire net_820;
wire net_821;
wire net_822;
wire net_823;
wire net_824;
wire net_825;
wire net_826;
wire net_828;
wire net_829;
wire net_830;
wire net_832;
wire net_833;
wire net_834;
wire net_835;
wire net_836;
wire net_837;
wire net_839;
wire net_840;
wire net_841;
wire net_843;
wire net_844;
wire net_845;
wire net_846;
wire net_847;
wire net_848;
wire net_849;
wire net_850;
wire net_851;
wire net_852;
wire net_853;
wire net_854;
wire net_856;
wire net_857;
wire net_858;
wire net_860;
wire net_861;
wire net_862;
wire net_863;
wire net_864;
wire net_865;
wire net_867;
wire net_868;
wire net_869;
wire net_871;
wire net_872;
wire net_873;
wire net_874;
wire net_875;
wire net_876;
wire net_877;
wire net_878;
wire net_879;
wire net_881;
wire net_882;
wire net_883;
wire net_885;
wire net_886;
wire net_887;
wire net_888;
wire net_889;
wire net_890;
wire net_892;
wire net_893;
wire net_894;
wire net_896;
wire net_897;
wire net_898;
wire net_899;
wire net_900;
wire net_901;
wire net_902;
wire net_903;
wire net_904;
wire net_906;
wire net_907;
wire nc16129;
wire nc16130;
wire nc16131;
wire nc16132;
wire nc16133;
wire nc16134;
wire nc16135;
wire nc16136;
wire nc16137;
wire nc16138;
wire nc16139;
wire nc16140;
wire nc16141;
wire nc16142;
wire nc16143;
wire nc16144;
wire nc16145;
wire nc16146;
wire nc16147;
wire nc16148;
wire nc16149;
wire nc16150;
wire nc16151;
wire nc16152;
wire nc16153;
wire nc16154;
wire nc16155;
wire nc16156;
wire nc16157;
wire nc16158;
wire nc16159;
wire nc16160;
wire nc16161;
wire nc16162;
wire nc16163;
wire nc16164;
wire nc16165;
wire nc16166;
wire nc16167;
wire nc16168;
wire nc16169;
wire nc16170;
wire nc16171;
wire nc16172;
wire nc16173;
wire nc16174;
wire nc16175;
wire nc16176;
wire nc16177;
wire nc16178;
wire nc16179;
wire nc16180;
wire nc16181;
wire nc16182;
wire nc16183;
wire nc16184;
wire nc16185;
wire nc16186;
wire nc16187;
wire nc16188;
wire nc16189;
wire nc16190;
wire nc16191;
wire nc16192;
wire nc16193;
wire nc16194;
wire nc16195;
wire nc16196;
wire nc16197;
wire nc16198;
wire nc16199;
wire nc16200;
wire nc16201;
wire nc16202;
wire nc16203;
wire nc16204;
wire nc16205;
wire nc16206;
wire nc16207;
wire nc16208;
wire nc16209;
wire nc16210;
wire nc16211;
wire nc16212;
wire nc16213;
wire nc16214;
wire nc16215;
wire nc16216;
wire nc16217;
wire nc16218;
wire nc16219;
wire nc16220;
wire nc16221;
wire nc16222;
wire nc16223;
wire nc16224;
wire nc16225;
wire nc16226;
wire nc16227;
wire nc16228;
wire nc16229;
wire nc16230;
wire nc16231;
wire nc16232;
wire nc16233;
wire nc16234;
wire nc16235;
wire nc16236;
wire nc16237;
wire nc16238;
wire nc16239;
wire nc16240;
wire nc16241;
wire nc16242;
wire nc16243;
wire nc16244;
wire nc16245;
wire nc16246;
wire nc16247;
wire nc16248;
wire nc16249;
wire nc16250;
wire nc16251;
wire nc16252;
wire nc16253;
wire nc16254;
wire nc16255;
wire nc16256;
wire nc16257;
wire nc16258;
wire nc16259;
wire nc16260;
wire nc16261;
wire nc16262;
wire nc16263;
wire nc16264;
wire nc16265;
wire nc16266;
wire nc16267;
wire nc16268;
wire nc16269;
wire nc16270;
wire nc16271;
wire nc16272;
wire nc16273;
wire nc16274;
wire nc16275;
wire nc16276;
wire nc16277;
wire nc16278;
wire nc16279;
wire nc16280;
wire nc16281;
wire nc16282;
wire nc16283;
wire nc16284;
wire nc16285;
wire nc16286;
wire nc16287;
wire nc16288;
wire nc16289;
wire nc16290;
wire nc16291;
wire nc16292;
wire nc16293;
wire nc16294;
wire nc16295;
wire nc16296;
wire nc16297;
wire nc16298;
wire nc16299;
wire nc16300;
wire nc16301;
wire nc16302;
wire nc16303;
wire nc16304;
wire nc16305;
wire nc16306;
wire nc16307;
wire nc16308;
wire nc16309;
wire nc16310;
wire nc16311;
wire nc16312;
wire nc16313;
wire nc16314;
wire nc16315;
wire nc16316;
wire nc16317;
wire nc16318;
wire nc16319;
wire nc16320;
wire nc16321;
wire nc16322;
wire nc16323;
wire nc16324;
wire nc16325;
wire nc16326;
wire nc16327;
wire nc16328;
wire nc16329;
wire nc16330;
wire nc16331;
wire nc16332;
wire nc16333;
wire nc16334;
wire nc16335;
wire nc16336;
wire nc16337;
wire nc16338;
wire nc16339;
wire nc16340;
wire nc16341;
wire nc16342;
wire nc16343;
wire nc16344;
wire nc16345;
wire nc16346;
wire nc16347;
wire nc16348;
wire nc16349;
wire nc16350;
wire nc16351;
wire nc16352;
wire nc16353;
wire nc16354;
wire nc16355;
wire nc16356;
wire nc16357;
wire nc16358;
wire nc16359;
wire nc16360;
wire nc16361;
wire nc16362;
wire nc16363;
wire nc16364;
wire nc16365;
wire nc16366;
wire nc16367;
wire nc16368;
wire nc16369;
wire nc16370;
wire nc16371;
wire nc16372;
wire nc16373;
wire nc16374;
wire nc16375;
wire nc16376;
wire nc16377;
wire nc16378;
wire nc16379;
wire nc16380;
wire nc16381;
wire nc16382;
wire nc16383;
wire nc16384;
wire nc16385;
wire nc16386;
wire nc16387;
wire nc16388;
wire nc16389;
wire nc16390;
wire nc16391;
wire nc16392;
wire nc16393;
wire nc16394;
wire nc16395;
wire nc16396;
wire nc16397;
wire nc16398;
wire nc16399;
wire nc16400;
wire nc16401;
wire nc16402;
wire nc16403;
wire nc16404;
wire nc16405;
wire nc16406;
wire nc16407;
wire nc16408;
wire nc16409;
wire nc16410;
wire nc16411;
wire nc16412;
wire nc16413;
wire nc16414;
wire nc16415;
wire nc16416;
wire nc16417;
wire nc16418;
wire nc16419;
wire nc16420;
wire nc16421;
wire nc16422;
wire nc16423;
wire nc16424;
wire nc16425;
wire nc16426;
wire nc16427;
wire nc16428;
wire nc16429;
wire nc16430;
wire nc16431;
wire nc16432;
wire nc16433;
wire nc16434;
wire nc16435;
wire nc16436;
wire nc16437;
wire nc16438;
wire nc16439;
wire nc16440;
wire nc16441;
wire nc16442;
wire nc16443;
wire nc16444;
wire nc16445;
wire nc16446;
wire nc16447;
wire nc16448;
wire nc16449;
wire nc16450;
wire nc16451;
wire nc16452;
wire nc16453;
wire nc16454;
wire nc16455;
wire nc16456;
wire nc16457;
wire nc16458;
wire nc16459;
wire nc16460;
wire nc16461;
wire nc16462;
wire nc16463;
wire nc16464;
wire nc16465;
wire nc16466;
wire nc16467;
wire nc16468;
wire nc16469;
wire nc16470;
wire nc16471;
wire nc16472;
wire nc16473;
wire nc16474;
wire nc16475;
wire nc16476;
wire nc16477;
wire nc16478;
wire nc16479;
wire nc16480;
wire nc16481;
wire nc16482;
wire nc16483;
wire nc16484;
wire nc16485;
wire nc16486;
wire nc16487;
wire nc16488;
wire nc16489;
wire nc16490;
wire nc16491;
wire nc16492;
wire nc16493;
wire nc16494;
wire nc16495;
wire nc16496;
wire nc16497;
wire nc16498;
wire nc16499;
wire nc16500;
wire nc16501;
wire nc16502;
wire nc16503;
wire nc16504;
wire nc16505;
wire nc16506;
wire nc16507;
wire nc16508;
wire nc16509;
wire nc16510;
wire nc16511;
wire nc16512;
wire nc16513;
wire nc16514;
wire nc16515;
wire nc16516;
wire nc16517;
wire nc16518;
wire nc16519;
wire nc16520;
wire nc16521;
wire nc16522;
wire nc16523;
wire nc16524;
wire nc16525;
wire nc16526;
wire nc16527;
wire nc16528;
wire nc16529;
wire nc16530;
wire nc16531;
wire nc16532;
wire nc16533;
wire nc16534;
wire nc16535;
wire nc16536;
wire nc16537;
wire nc16538;
wire nc16539;
wire nc16540;
wire nc16541;
wire nc16542;
wire nc16543;
wire nc16544;
wire nc16545;
wire nc16546;
wire nc16547;
wire nc16548;
wire nc16549;
wire nc16550;
wire nc16551;
wire nc16552;
wire nc16553;
wire nc16554;
wire nc16555;
wire nc16556;
wire nc16557;
wire nc16558;
wire nc16559;
wire nc16560;
wire nc16561;
wire nc16562;
wire nc16563;
wire nc16564;
wire nc16565;
wire nc16566;
wire nc16567;
wire nc16568;
wire nc16569;
wire nc16570;
wire nc16571;
wire nc16572;
wire nc16573;
wire nc16574;
wire nc16575;
wire nc16576;
wire nc16577;
wire nc16578;
wire nc16579;
wire nc16580;
wire nc16581;
wire nc16582;
wire nc16583;
wire nc16584;
wire nc16585;
wire nc16586;
wire nc16587;
wire nc16588;
wire nc16589;
wire nc16590;
wire nc16591;
wire nc16592;
wire nc16593;
wire nc16594;
wire nc16595;
wire nc16596;
wire nc16597;
wire nc16598;
wire nc16599;
wire nc16600;
wire nc16601;
wire nc16602;
wire nc16603;
wire nc16604;
wire nc16605;
wire nc16606;
wire nc16607;
wire nc16608;
wire nc16609;
wire nc16610;
wire nc16611;
wire nc16612;
wire nc16613;
wire nc16614;
wire nc16615;
wire nc16616;
wire nc16617;
wire nc16618;
wire nc16619;
wire nc16620;
wire nc16621;
wire nc16622;
wire nc16623;
wire nc16624;
wire nc16625;
wire nc16626;
wire nc16627;
wire nc16628;
wire nc16629;
wire nc16630;
wire nc16631;
wire nc16632;
wire nc16633;
wire nc16634;
wire nc16635;
wire nc16636;
wire nc16637;
wire nc16638;
wire nc16639;
wire nc16640;
wire nc16641;
wire nc16642;
wire nc16643;
wire nc16644;
wire nc16645;
wire nc16646;
wire nc16647;
wire nc16648;
wire nc16649;
wire nc16650;
wire nc16651;
wire nc16652;
wire nc16653;
wire nc16654;
wire nc16655;
wire nc16656;
wire nc16657;
wire nc16658;
wire nc16659;
wire nc16660;
wire nc16661;
wire nc16662;
wire nc16663;
wire nc16664;
wire nc16665;
wire nc16666;
wire nc16667;
wire nc16668;
wire nc16669;
wire nc16670;
wire nc16671;
wire nc16672;
wire nc16673;
wire nc16674;
wire nc16675;
wire nc16676;
wire nc16677;
wire nc16678;
wire nc16679;
wire nc16680;
wire nc16681;
wire nc16682;
wire nc16683;
wire nc16684;
wire nc16685;
wire nc16686;
wire nc16687;
wire nc16688;
wire nc16689;
wire nc16690;
wire nc16691;
wire nc16692;
wire nc16693;
wire nc16694;
wire nc16695;
wire nc16696;
wire nc16697;
wire nc16698;
wire nc16699;
wire nc16700;
wire nc16701;
wire nc16702;
wire nc16703;
wire nc16704;
wire nc16705;
wire nc16706;
wire nc16707;
wire nc16708;
wire nc16709;
wire nc16710;
wire nc16711;
wire nc16712;
wire nc16713;
wire nc16714;
wire nc16715;
wire nc16716;
wire nc16717;
wire nc16718;
wire nc16719;
wire nc16720;
wire nc16721;
wire nc16722;
wire nc16723;
wire nc16724;
wire nc16725;
wire nc16726;
wire nc16727;
wire nc16728;
wire nc16729;
wire nc16730;
wire nc16731;
wire nc16732;
wire nc16733;
wire nc16734;
wire nc16735;
wire nc16736;
wire nc16737;
wire nc16738;
wire nc16739;
wire nc16740;
wire nc16741;
wire nc16742;
wire nc16743;
wire nc16744;
wire nc16745;
wire nc16746;
wire nc16747;
wire nc16748;
wire nc16749;
wire nc16750;
wire nc16751;
wire nc16752;
wire nc16753;
wire nc16754;
wire nc16755;
wire nc16756;
wire nc16757;
wire nc16758;
wire nc16759;
wire nc16760;
wire nc16761;
wire nc16762;
wire nc16763;
wire nc16764;
wire nc16765;
wire nc16766;
wire nc16767;
wire nc16768;
wire nc16769;
wire nc16770;
wire nc16771;
wire nc16772;
wire nc16773;
wire nc16774;
wire nc16775;
wire nc16776;
wire nc16777;
wire nc16778;
wire nc16779;
wire nc16780;
wire nc16781;
wire nc16782;
wire nc16783;
wire nc16784;
wire nc16785;
wire nc16786;
wire nc16787;
wire nc16788;
wire nc16789;
wire nc16790;
wire nc16791;
wire nc16792;
wire nc16793;
wire nc16794;
wire nc16795;
wire nc16796;
wire nc16797;
wire nc16798;
wire nc16799;
wire nc16800;
wire nc16801;
wire nc16802;
wire nc16803;
wire nc16804;
wire nc16805;
wire nc16806;
wire nc16807;
wire nc16808;
wire nc16809;
wire nc16810;
wire nc16811;
wire nc16812;
wire nc16813;
wire nc16814;
wire nc16815;
wire nc16816;
wire nc16817;
wire nc16818;
wire nc16819;
wire nc16820;
wire nc16821;
wire nc16822;
wire nc16823;
wire nc16824;
wire nc16825;
wire nc16826;
wire nc16827;
wire nc16828;
wire nc16829;
wire nc16830;
wire nc16831;
wire nc16832;
wire nc16833;
wire nc16834;
wire nc16835;
wire nc16836;
wire nc16837;
wire nc16838;
wire nc16839;
wire nc16840;
wire nc16841;
wire nc16842;
wire nc16843;
wire nc16844;
wire nc16845;
wire nc16846;
wire nc16847;
wire nc16848;
wire nc16849;
wire nc16850;
wire nc16851;
wire nc16852;
wire nc16853;
wire nc16854;
wire nc16855;
wire nc16856;
wire nc16857;
wire nc16858;
wire nc16859;
wire nc16860;
wire nc16861;
wire nc16862;
wire nc16863;
wire nc16864;
wire nc16865;
wire nc16866;
wire nc16867;
wire nc16868;
wire nc16869;
wire nc16870;
wire nc16871;
wire nc16872;
wire nc16873;
wire nc16874;
wire nc16875;
wire nc16876;
wire nc16877;
wire nc16878;
wire nc16879;
wire nc16880;
wire nc16881;
wire nc16882;
wire nc16883;
wire nc16884;
wire nc16885;
wire nc16886;
wire nc16887;
wire nc16888;
wire nc16889;
wire nc16890;
wire nc16891;
wire nc16892;
wire nc16893;
wire nc16894;
wire nc16895;
wire nc16896;
wire nc16897;
wire nc16898;
wire nc16899;
wire nc16900;
wire nc16901;
wire nc16902;
wire nc16903;
wire nc16904;
wire nc16905;
wire nc16906;
wire nc16907;
wire nc16908;
wire nc16909;
wire nc16910;
wire nc16911;
wire nc16912;
wire nc16913;
wire nc16914;
wire nc16915;
wire nc16916;
wire nc16917;
wire nc16918;
wire nc16919;
wire nc16920;
wire nc16921;
wire nc16922;
wire nc16923;
wire nc16924;
wire nc16925;
wire nc16926;
wire nc16927;
wire nc16928;
wire nc16929;
wire nc16930;
wire nc16931;
wire nc16932;
wire nc16933;
wire nc16934;
wire nc16935;
wire nc16936;
wire nc16937;
wire nc16938;
wire nc16939;
wire nc16940;
wire nc16941;
wire nc16942;
wire nc16943;
wire nc16944;
wire nc16945;
wire nc16946;
wire nc16947;
wire nc16948;
wire nc16949;
wire nc16950;
wire nc16951;
wire nc16952;
wire nc16953;
wire nc16954;
wire nc16955;
wire nc16956;
wire nc16957;
wire nc16958;
wire nc16959;
wire nc16960;
wire nc16961;
wire nc16962;
wire nc16963;
wire nc16964;
wire nc16965;
wire nc16966;
wire nc16967;
wire nc16968;
wire nc16969;
wire nc16970;
wire nc16971;
wire nc16972;
wire nc16973;
wire nc16974;
wire nc16975;
wire nc16976;
wire nc16977;
wire nc16978;
wire nc16979;
wire nc16980;
wire nc16981;
wire nc16982;
wire nc16983;
wire nc16984;
wire nc16985;
wire nc16986;
wire nc16987;
wire nc16988;
wire nc16989;
wire nc16990;
wire nc16991;
wire nc16992;
wire nc16993;
wire nc16994;
wire nc16995;
wire nc16996;
wire nc16997;
wire nc16998;
wire nc16999;
wire nc17000;
wire nc17001;
wire nc17002;
wire nc17003;
wire nc17004;
wire nc17005;
wire nc17006;
wire nc17007;
wire nc17008;
wire nc17009;
wire nc17010;
wire nc17011;
wire nc17012;
wire nc17013;
wire nc17014;
wire nc17015;
wire nc17016;
wire nc17017;
wire nc17018;
wire nc17019;
wire nc17020;
wire nc17021;
wire nc17022;
wire nc17023;
wire nc17024;
wire nc17025;
wire nc17026;
wire nc17027;
wire nc17028;
wire nc17029;
wire nc17030;
wire nc17031;
wire nc17032;
wire nc17033;
wire nc17034;
wire nc17035;
wire nc17036;
wire nc17037;
wire nc17038;
wire nc17039;
wire nc17040;
wire nc17041;
wire nc17042;
wire nc17043;
wire nc17044;
wire nc17045;
wire nc17046;
wire nc17047;
wire nc17048;
wire nc17049;
wire nc17050;
wire nc17051;
wire nc17052;
wire nc17053;
wire nc17054;
wire nc17055;
wire nc17056;
wire nc17057;
wire nc17058;
wire nc17059;
wire nc17060;
wire nc17061;
wire nc17062;
wire nc17063;
wire nc17064;
wire nc17065;
wire nc17066;
wire nc17067;
wire nc17068;
wire nc17069;
wire nc17070;
wire nc17071;
wire nc17072;
wire nc17073;
wire nc17074;
wire nc17075;
wire nc17076;
wire nc17077;
wire nc17078;
wire nc17079;
wire nc17080;
wire nc17081;
wire nc17082;
wire nc17083;
wire nc17084;
wire nc17085;
wire nc17086;
wire nc17087;
wire nc17088;
wire nc17089;
wire nc17090;
wire nc17091;
wire nc17092;
wire nc17093;
wire nc17094;
wire nc17095;
wire nc17096;
wire nc17097;
wire nc17098;
wire nc17099;
wire nc17100;
wire nc17101;
wire nc17102;
wire nc17103;
wire nc17104;
wire nc17105;
wire nc17106;
wire nc17107;
wire nc17108;
wire nc17109;
wire nc17110;
wire nc17111;
wire nc17112;
wire nc17113;
wire nc17114;
wire nc17115;
wire nc17116;
wire nc17117;
wire nc17118;
wire nc17119;
wire nc17120;
wire nc17121;
wire nc17122;
wire nc17123;
wire nc17124;
wire nc17125;
wire nc17126;
wire nc17127;
wire nc17128;
wire nc17129;
wire nc17130;
wire nc17131;
wire nc17132;
wire nc17133;
wire nc17134;
wire nc17135;
wire nc17136;
wire nc17137;
wire nc17138;
wire nc17139;
wire nc17140;
wire nc17141;
wire nc17142;
wire nc17143;
wire nc17144;
wire nc17145;
wire nc17146;
wire nc17147;
wire nc17148;
wire nc17149;
wire nc17150;
wire nc17151;
wire nc17152;
wire nc17153;
wire nc17154;
wire nc17155;
wire nc17156;
wire nc17157;
wire nc17158;
wire nc17159;
wire nc17160;
wire nc17161;
wire nc17162;
wire nc17163;
wire nc17164;
wire nc17165;
wire nc17166;
wire nc17167;
wire nc17168;
wire nc17169;
wire nc17170;
wire nc17171;
wire nc17172;
wire nc17173;
wire nc17174;
wire nc17175;
wire nc17176;
wire nc17177;
wire nc17178;
wire nc17179;
wire nc17180;
wire nc17181;
wire nc17182;
wire nc17183;
wire nc17184;
wire nc17185;
wire nc17186;
wire nc17187;
wire nc17188;
wire nc17189;
wire nc17190;
wire nc17191;
wire nc17192;
wire nc17193;
wire nc17194;
wire nc17195;
wire nc17196;
wire nc17197;
wire nc17198;
wire nc17199;
wire nc17200;
wire nc17201;
wire nc17202;
wire nc17203;
wire nc17204;
wire nc17205;
wire nc17206;
wire nc17207;
wire nc17208;
wire nc17209;
wire nc17210;
wire nc17211;
wire nc17212;
wire nc17213;
wire nc17214;
wire nc17215;
wire nc17216;
wire nc17217;
wire nc17218;
wire nc17219;
wire nc17220;
wire nc17221;
wire nc17222;
wire nc17223;
wire nc17224;
wire nc17225;
wire nc17226;
wire nc17227;
wire nc17228;
wire nc17229;
wire nc17230;
wire nc17231;
wire nc17232;
wire nc17233;
wire nc17234;
wire nc17235;
wire nc17236;
wire nc17237;
wire nc17238;
wire nc17239;
wire nc17240;
wire nc17241;
wire nc17242;
wire nc17243;
wire nc17244;
wire nc17245;
wire nc17246;
wire nc17247;
wire nc17248;
wire nc17249;
wire nc17250;
wire nc17251;
wire nc17252;
wire nc17253;
wire nc17254;
wire nc17255;
wire nc17256;
wire nc17257;
wire nc17258;
wire nc17259;
wire nc17260;
wire nc17261;
wire nc17262;
wire nc17263;
wire nc17264;
wire nc17265;
wire nc17266;
wire nc17267;
wire nc17268;
wire nc17269;
wire nc17270;
wire nc17271;
wire nc17272;
wire nc17273;
wire nc17274;
wire nc17275;
wire nc17276;
wire nc17277;
wire nc17278;
wire nc17279;
wire nc17280;
wire nc17281;
wire nc17282;
wire nc17283;
wire nc17284;
wire nc17285;
wire nc17286;
wire nc17287;
wire nc17288;
wire nc17289;
wire nc17290;
wire nc17291;
wire nc17292;
wire nc17293;
wire nc17294;
wire nc17295;
wire nc17296;
wire nc17297;
wire nc17298;
wire nc17299;
wire nc17300;
wire nc17301;
wire nc17302;
wire nc17303;
wire nc17304;
wire nc17305;
wire nc17306;
wire nc17307;
wire nc17308;
wire nc17309;
wire nc17310;
wire nc17311;
wire nc17312;
wire nc17313;
wire nc17314;
wire nc17315;
wire nc17316;
wire nc17317;
wire nc17318;
wire nc17319;
wire nc17320;
wire nc17321;
wire nc17322;
wire nc17323;
wire nc17324;
wire nc17325;
wire nc17326;
wire nc17327;
wire nc17328;
wire nc17329;
wire nc17330;
wire nc17331;
wire nc17332;
wire nc17333;
wire nc17334;
wire nc17335;
wire nc17336;
wire nc17337;
wire nc17338;
wire nc17339;
wire nc17340;
wire nc17341;
wire nc17342;
wire nc17343;
wire nc17344;
wire nc17345;
wire nc17346;
wire nc17347;
wire nc17348;
wire nc17349;
wire nc17350;
wire nc17351;
wire nc17352;
wire nc17353;
wire nc17354;
wire nc17355;
wire nc17356;
wire nc17357;
wire nc17358;
wire nc17359;
wire nc17360;
wire nc17361;
wire nc17362;
wire nc17363;
wire nc17364;
wire nc17365;
wire nc17366;
wire nc17367;
wire nc17368;
wire nc17369;
wire nc17370;
wire nc17371;
wire nc17372;
wire nc17373;
wire nc17374;
wire nc17375;
wire nc17376;
wire nc17377;
wire nc17378;
wire nc17379;
wire nc17380;
wire nc17381;
wire nc17382;
wire nc17383;
wire nc17384;
wire nc17385;
wire nc17386;
wire nc17387;
wire nc17388;
wire nc17389;
wire nc17390;
wire nc17391;
wire nc17392;
wire nc17393;
wire nc17394;
wire nc17395;
wire nc17396;
wire nc17397;
wire nc17398;
wire nc17399;
wire nc17400;
wire nc17401;
wire nc17402;
wire nc17403;
wire nc17404;
wire nc17405;
wire nc17406;
wire nc17407;
wire nc17408;
wire nc17409;
wire nc17410;
wire nc17411;
wire nc17412;
wire nc17413;
wire nc17414;
wire nc17415;
wire nc17416;
wire nc17417;
wire nc17418;
wire nc17419;
wire nc17420;
wire nc17421;
wire nc17422;
wire nc17423;
wire nc17424;
wire nc17425;
wire nc17426;
wire nc17427;
wire nc17428;
wire nc17429;
wire nc17430;
wire nc17431;
wire nc17432;
wire nc17433;
wire nc17434;
wire nc17435;
wire nc17436;
wire nc17437;
wire nc17438;
wire nc17439;
wire nc17440;
wire nc17441;
wire nc17442;
wire nc17443;
wire nc17444;
wire nc17445;
wire nc17446;
wire nc17447;
wire nc17448;
wire nc17449;
wire nc17450;
wire nc17451;
wire nc17452;
wire nc17453;
wire nc17454;
wire nc17455;
wire nc17456;
wire nc17457;
wire nc17458;
wire nc17459;
wire nc17460;
wire nc17461;
wire nc17462;
wire nc17463;
wire nc17464;
wire nc17465;
wire nc17466;
wire nc17467;
wire nc17468;
wire nc17469;
wire nc17470;
wire nc17471;
wire nc17472;
wire nc17473;
wire nc17474;
wire nc17475;
wire nc17476;
wire nc17477;
wire nc17478;
wire nc17479;
wire nc17480;
wire nc17481;
wire nc17482;
wire nc17483;
wire nc17484;
wire nc17485;
wire nc17486;
wire nc17487;
wire nc17488;
wire nc17489;
wire nc17490;
wire nc17491;
wire nc17492;
wire nc17493;
wire nc17494;
wire nc17495;
wire nc17496;
wire nc17497;
wire nc17498;
wire nc17499;
wire nc17500;
wire nc17501;
wire nc17502;
wire nc17503;
wire nc17504;
wire nc17505;
wire nc17506;
wire nc17507;
wire nc17508;
wire nc17509;
wire nc17510;
wire nc17511;
wire nc17512;
wire nc17513;
wire nc17514;
wire nc17515;
wire nc17516;
wire nc17517;
wire nc17518;
wire nc17519;
wire nc17520;
wire nc17521;
wire nc17522;
wire nc17523;
wire nc17524;
wire nc17525;
wire nc17526;
wire nc17527;
wire nc17528;
wire nc17529;
wire nc17530;
wire nc17531;
wire nc17532;
wire nc17533;
wire nc17534;
wire nc17535;
wire nc17536;
wire nc17537;
wire nc17538;
wire nc17539;
wire nc17540;
wire nc17541;
wire nc17542;
wire nc17543;
wire nc17544;
wire nc17545;
wire nc17546;
wire nc17547;
wire nc17548;
wire nc17549;
wire nc17550;
wire nc17551;
wire nc17552;
wire nc17553;
wire nc17554;
wire nc17555;
wire nc17556;
wire nc17557;
wire nc17558;
wire nc17559;
wire nc17560;
wire nc17561;
wire nc17562;
wire nc17563;
wire nc17564;
wire nc17565;
wire nc17566;
wire nc17567;
wire nc17568;
wire nc17569;
wire nc17570;
wire nc17571;
wire nc17572;
wire nc17573;
wire nc17574;
wire nc17575;
wire nc17576;
wire nc17577;
wire nc17578;
wire nc17579;
wire nc17580;
wire nc17581;
wire nc17582;
wire nc17583;
wire nc17584;
wire nc17585;
wire nc17586;
wire nc17587;
wire nc17588;
wire nc17589;
wire nc17590;
wire nc17591;
wire nc17592;
wire nc17593;
wire nc17594;
wire nc17595;
wire nc17596;
wire nc17597;
wire nc17598;
wire nc17599;
wire nc17600;
wire nc17601;
wire nc17602;
wire nc17603;
wire nc17604;
wire nc17605;
wire nc17606;
wire nc17607;
wire nc17608;
wire nc17609;
wire nc17610;
wire nc17611;
wire nc17612;
wire nc17613;
wire nc17614;
wire nc17615;
wire nc17616;
wire nc17617;
wire nc17618;
wire nc17619;
wire nc17620;
wire nc17621;
wire nc17622;
wire nc17623;
wire nc17624;
wire nc17625;
wire nc17626;
wire nc17627;
wire nc17628;
wire nc17629;
wire nc17630;
wire nc17631;
wire nc17632;
wire nc17633;
wire nc17634;
wire nc17635;
wire nc17636;
wire nc17637;
wire nc17638;
wire nc17639;
wire nc17640;
wire nc17641;
wire nc17642;
wire nc17643;
wire nc17644;
wire nc17645;
wire nc17646;
wire nc17647;
wire nc17648;
wire nc17649;
wire nc17650;
wire nc17651;
wire nc17652;
wire nc17653;
wire nc17654;
wire nc17655;
wire nc17656;
wire nc17657;
wire nc17658;
wire nc17659;
wire nc17660;
wire nc17661;
wire nc17662;
wire nc17663;
wire nc17664;
wire nc17665;
wire nc17666;
wire nc17667;
wire nc17668;
wire nc17669;
wire nc17670;
wire nc17671;
wire nc17672;
wire nc17673;
wire nc17674;
wire nc17675;
wire nc17676;
wire nc17677;
wire nc17678;
wire nc17679;
wire nc17680;
wire nc17681;
wire nc17682;
wire nc17683;
wire nc17684;
wire nc17685;
wire nc17686;
wire nc17687;
wire nc17688;
wire nc17689;
wire nc17690;
wire nc17691;
wire nc17692;
wire nc17693;
wire nc17694;
wire nc17695;
wire nc17696;
wire nc17697;
wire nc17698;
wire nc17699;
wire nc17700;
wire nc17701;
wire nc17702;
wire nc17703;
wire nc17704;
wire nc17705;
wire nc17706;
wire nc17707;
wire nc17708;
wire nc17709;
wire nc17710;
wire nc17711;
wire nc17712;
wire nc17713;
wire nc17714;
wire nc17715;
wire nc17716;
wire nc17717;
wire nc17718;
wire nc17719;
wire nc17720;
wire nc17721;
wire nc17722;
wire nc17723;
wire nc17724;
wire nc17725;
wire nc17726;
wire nc17727;
wire nc17728;
wire nc17729;
wire nc17730;
wire nc17731;
wire nc17732;
wire nc17733;
wire nc17734;
wire nc17735;
wire nc17736;
wire nc17737;
wire nc17738;
wire nc17739;
wire nc17740;
wire nc17741;
wire nc17742;
wire nc17743;
wire nc17744;
wire nc17745;
wire nc17746;
wire nc17747;
wire nc17748;
wire nc17749;
wire nc17750;
wire nc17751;
wire nc17752;
wire nc17753;
wire nc17754;
wire nc17755;
wire nc17756;
wire nc17757;
wire nc17758;
wire nc17759;
wire nc17760;
wire nc17761;
wire nc17762;
wire nc17763;
wire nc17764;
wire nc17765;
wire nc17766;
wire nc17767;
wire nc17768;
wire nc17769;
wire nc17770;
wire nc17771;
wire nc17772;
wire nc17773;
wire nc17774;
wire nc17775;
wire nc17776;
wire nc17777;
wire nc17778;
wire nc17779;
wire nc17780;
wire nc17781;
wire nc17782;
wire nc17783;
wire nc17784;
wire nc17785;
wire nc17786;
wire nc17787;
wire nc17788;
wire nc17789;
wire nc17790;
wire nc17791;
wire nc17792;
wire nc17793;
wire nc17794;
wire nc17795;
wire nc17796;
wire nc17797;
wire nc17798;
wire nc17799;
wire nc17800;
wire nc17801;
wire nc17802;
wire nc17803;
wire nc17804;
wire nc17805;
wire nc17806;
wire nc17807;
wire nc17808;
wire nc17809;
wire nc17810;
wire nc17811;
wire nc17812;
wire nc17813;
wire nc17814;
wire nc17815;
wire nc17816;
wire nc17817;
wire nc17818;
wire nc17819;
wire nc17820;
wire nc17821;
wire nc17822;
wire nc17823;
wire nc17824;
wire nc17825;
wire nc17826;
wire nc17827;
wire nc17828;
wire nc17829;
wire nc17830;
wire nc17831;
wire nc17832;
wire nc17833;
wire nc17834;
wire nc17835;
wire nc17836;
wire nc17837;
wire nc17838;
wire nc17839;
wire nc17840;
wire nc17841;
wire nc17842;
wire nc17843;
wire nc17844;
wire nc17845;
wire nc17846;
wire nc17847;
wire nc17848;
wire nc17849;
wire nc17850;
wire nc17851;
wire nc17852;
wire nc17853;
wire nc17854;
wire nc17855;
wire nc17856;
wire nc17857;
wire nc17858;
wire nc17859;
wire nc17860;
wire nc17861;
wire nc17862;
wire nc17863;
wire nc17864;
wire nc17865;
wire nc17866;
wire nc17867;
wire nc17868;
wire nc17869;
wire nc17870;
wire nc17871;
wire nc17872;
wire nc17873;
wire nc17874;
wire nc17875;
wire nc17876;
wire nc17877;
wire nc17878;
wire nc17879;
wire nc17880;
wire nc17881;
wire nc17882;
wire nc17883;
wire nc17884;
wire nc17885;
wire nc17886;
wire nc17887;
wire nc17888;
wire nc17889;
wire nc17890;
wire nc17891;
wire nc17892;
wire nc17893;
wire nc17894;
wire nc17895;
wire nc17896;
wire nc17897;
wire nc17898;
wire nc17899;
wire nc17900;
wire nc17901;
wire nc17902;
wire nc17903;
wire nc17904;
wire nc17905;
wire nc17906;
wire nc17907;
wire nc17908;
wire nc17909;
wire nc17910;
wire nc17911;
wire nc17912;
wire nc17913;
wire nc17914;
wire nc17915;
wire nc17916;
wire nc17917;
wire nc17918;
wire nc17919;
wire nc17920;
wire nc17921;
wire nc17922;
wire nc17923;
wire nc17924;
wire nc17925;
wire nc17926;
wire nc17927;
wire nc17928;
wire nc17929;
wire nc17930;
wire nc17931;
wire nc17932;
wire nc17933;
wire nc17934;
wire nc17935;
wire nc17936;
wire nc17937;
wire nc17938;
wire nc17939;
wire nc17940;
wire nc17941;
wire nc17942;
wire nc17943;
wire nc17944;
wire nc17945;
wire nc17946;
wire nc17947;
wire nc17948;
wire nc17949;
wire nc17950;
wire nc17951;
wire nc17952;
wire nc17953;
wire nc17954;
wire nc17955;
wire nc17956;
wire nc17957;
wire nc17958;
wire nc17959;
wire nc17960;
wire nc17961;
wire nc17962;
wire nc17963;
wire nc17964;
wire nc17965;
wire nc17966;
wire nc17967;
wire nc17968;
wire nc17969;
wire nc17970;
wire nc17971;
wire nc17972;
wire nc17973;
wire nc17974;
wire nc17975;
wire nc17976;
wire nc17977;
wire nc17978;
wire nc17979;
wire nc17980;
wire nc17981;
wire nc17982;
wire nc17983;
wire nc17984;
wire nc17985;
wire nc17986;
wire nc17987;
wire nc17988;
wire nc17989;
wire nc17990;
wire nc17991;
wire nc17992;
wire nc17993;
wire nc17994;
wire nc17995;
wire nc17996;
wire nc17997;
wire nc17998;
wire nc17999;
wire nc18000;
wire nc18001;
wire nc18002;
wire nc18003;
wire nc18004;
wire nc18005;
wire nc18006;
wire nc18007;
wire nc18008;
wire nc18009;
wire nc18010;
wire nc18011;
wire nc18012;
wire nc18013;
wire nc18014;
wire nc18015;
wire nc18016;
wire nc18017;
wire nc18018;
wire nc18019;
wire nc18020;
wire nc18021;
wire nc18022;
wire nc18023;
wire nc18024;
wire nc18025;
wire nc18026;
wire nc18027;
wire nc18028;
wire nc18029;
wire nc18030;
wire nc18031;
wire nc18032;
wire nc18033;
wire nc18034;
wire nc18035;
wire nc18036;
wire nc18037;
wire nc18038;
wire nc18039;
wire nc18040;
wire nc18041;
wire nc18042;
wire nc18043;
wire nc18044;
wire nc18045;
wire nc18046;
wire nc18047;
wire nc18048;
wire nc18049;
wire nc18050;
wire nc18051;
wire nc18052;
wire nc18053;
wire nc18054;
wire nc18055;
wire nc18056;
wire nc18057;
wire nc18058;
wire nc18059;
wire nc18060;
wire nc18061;
wire nc18062;
wire nc18063;
wire nc18064;
wire nc18065;
wire nc18066;
wire nc18067;
wire nc18068;
wire nc18069;
wire nc18070;
wire nc18071;
wire nc18072;
wire nc18073;
wire nc18074;
wire nc18075;
wire nc18076;
wire nc18077;
wire nc18078;
wire nc18079;
wire nc18080;
wire nc18081;
wire nc18082;
wire nc18083;
wire nc18084;
wire nc18085;
wire nc18086;
wire nc18087;
wire nc18088;
wire nc18089;
wire nc18090;
wire nc18091;
wire nc18092;
wire nc18093;
wire nc18094;
wire nc18095;
wire nc18096;
wire nc18097;
wire nc18098;
wire nc18099;
wire nc18100;
wire nc18101;
wire nc18102;
wire nc18103;
wire nc18104;
wire nc18105;
wire nc18106;
wire nc18107;
wire nc18108;
wire nc18109;
wire nc18110;
wire nc18111;
wire nc18112;
wire nc18113;
wire nc18114;
wire nc18115;
wire nc18116;
wire nc18117;
wire nc18118;
wire nc18119;
wire nc18120;
wire nc18121;
wire nc18122;
wire nc18123;
wire nc18124;
wire nc18125;
wire nc18126;
wire nc18127;
wire nc18128;
wire nc18129;
wire nc18130;
wire nc18131;
wire nc18132;
wire nc18133;
wire nc18134;
wire nc18135;
wire nc18136;
wire nc18137;
wire nc18138;
wire nc18139;
wire nc18140;
wire nc18141;
wire nc18142;
wire nc18143;
wire nc18144;
wire nc18145;
wire nc18146;
wire nc18147;
wire nc18148;
wire nc18149;
wire nc18150;
wire nc18151;
wire nc18152;
wire nc18153;
wire nc18154;
wire nc18155;
wire nc18156;
wire nc18157;
wire nc18158;
wire nc18159;
wire nc18160;
wire nc18161;
wire nc18162;
wire nc18163;
wire nc18164;
wire nc18165;
wire nc18166;
wire nc18167;
wire nc18168;
wire nc18169;
wire nc18170;
wire nc18171;
wire nc18172;
wire nc18173;
wire nc18174;
wire nc18175;
wire nc18176;
wire nc18177;
wire nc18178;
wire nc18179;
wire nc18180;
wire nc18181;
wire nc18182;
wire nc18183;
wire nc18184;
wire nc18185;
wire nc18186;
wire nc18187;
wire nc18188;
wire nc18189;
wire nc18190;
wire nc18191;
wire nc18192;
wire nc18193;
wire nc18194;
wire nc18195;
wire nc18196;
wire nc18197;
wire nc18198;
wire nc18199;
wire nc18200;
wire nc18201;
wire nc18202;
wire nc18203;
wire nc18204;
wire nc18205;
wire nc18206;
wire nc18207;
wire nc18208;
wire nc18209;
wire nc18210;
wire nc18211;
wire nc18212;
wire nc18213;
wire nc18214;
wire nc18215;
wire nc18216;
wire nc18217;
wire nc18218;
wire nc18219;
wire nc18220;
wire nc18221;
wire nc18222;
wire nc18223;
wire nc18224;
wire nc18225;
wire nc18226;
wire nc18227;
wire nc18228;
wire nc18229;
wire nc18230;
wire nc18231;
wire nc18232;
wire nc18233;
wire nc18234;
wire nc18235;
wire nc18236;
wire nc18237;
wire nc18238;
wire nc18239;
wire nc18240;
wire nc18241;
wire nc18242;
wire nc18243;
wire nc18244;
wire nc18245;
wire nc18246;
wire nc18247;
wire nc18248;
wire nc18249;
wire nc18250;
wire nc18251;
wire nc18252;
wire nc18253;
wire nc18254;
wire nc18255;
wire nc18256;
wire nc18257;
wire nc18258;
wire nc18259;
wire nc18260;
wire nc18261;
wire nc18262;
wire nc18263;
wire nc18264;
wire nc18265;
wire nc18266;
wire nc18267;
wire nc18268;
wire nc18269;
wire nc18270;
wire nc18271;
wire nc18272;
wire nc18273;
wire nc18274;
wire nc18275;
wire nc18276;
wire nc18277;
wire nc18278;
wire nc18279;
wire nc18280;
wire nc18281;
wire nc18282;
wire nc18283;
wire nc18284;
wire nc18285;
wire nc18286;
wire nc18287;
wire nc18288;
wire nc18289;
wire nc18290;
wire nc18291;
wire nc18292;
wire nc18293;
wire nc18294;
wire nc18295;
wire nc18296;
wire nc18297;
wire nc18298;
wire nc18299;
wire nc18300;
wire nc18301;
wire nc18302;
wire nc18303;
wire nc18304;
wire nc18305;
wire nc18306;
wire nc18307;
wire nc18308;
wire nc18309;
wire nc18310;
wire nc18311;
wire nc18312;
wire nc18313;
wire nc18314;
wire nc18315;
wire nc18316;
wire nc18317;
wire nc18318;
wire nc18319;
wire nc18320;
wire nc18321;
wire nc18322;
wire nc18323;
wire nc18324;
wire nc18325;
wire nc18326;
wire nc18327;
wire nc18328;
wire nc18329;
wire nc18330;
wire nc18331;
wire nc18332;
wire nc18333;
wire nc18334;
wire nc18335;
wire nc18336;
wire nc18337;
wire nc18338;
wire nc18339;
wire nc18340;
wire nc18341;
wire nc18342;
wire nc18343;
wire nc18344;
wire nc18345;
wire nc18346;
wire nc18347;
wire nc18348;
wire nc18349;
wire nc18350;
wire nc18351;
wire nc18352;
wire nc18353;
wire nc18354;
wire nc18355;
wire nc18356;
wire nc18357;
wire nc18358;
wire nc18359;
wire nc18360;
wire nc18361;
wire nc18362;
wire nc18363;
wire nc18364;
wire nc18365;
wire nc18366;
wire nc18367;
wire nc18368;
wire nc18369;
wire nc18370;
wire nc18371;
wire nc18372;
wire nc18373;
wire nc18374;
wire nc18375;
wire nc18376;
wire nc18377;
wire nc18378;
wire nc18379;
wire nc18380;
wire nc18381;
wire nc18382;
wire nc18383;
wire nc18384;
wire nc18385;
wire nc18386;
wire nc18387;
wire nc18388;
wire nc18389;
wire nc18390;
wire nc18391;
wire nc18392;
wire nc18393;
wire nc18394;
wire nc18395;
wire nc18396;
wire nc18397;
wire nc18398;
wire nc18399;
wire nc18400;
wire nc18401;
wire nc18402;
wire nc18403;
wire nc18404;
wire nc18405;
wire nc18406;
wire nc18407;
wire nc18408;
wire nc18409;
wire nc18410;
wire nc18411;
wire nc18412;
wire nc18413;
wire nc18414;
wire nc18415;
wire nc18416;
wire nc18417;
wire nc18418;
wire nc18419;
wire nc18420;
wire nc18421;
wire nc18422;
wire nc18423;
wire nc18424;
wire nc18425;
wire nc18426;
wire nc18427;
wire nc18428;
wire nc18429;
wire nc18430;
wire nc18431;
wire nc18432;
wire nc18433;
wire nc18434;
wire nc18435;
wire nc18436;
wire nc18437;
wire nc18438;
wire nc18439;
wire nc18440;
wire nc18441;
wire nc18442;
wire nc18443;
wire nc18444;
wire nc18445;
wire nc18446;
wire nc18447;
wire nc18448;
wire nc18449;
wire nc18450;
wire nc18451;
wire nc18452;
wire nc18453;
wire nc18454;
wire nc18455;
wire nc18456;
wire nc18457;
wire nc18458;
wire nc18459;
wire nc18460;
wire nc18461;
wire nc18462;
wire nc18463;
wire nc18464;
wire nc18465;
wire nc18466;
wire nc18467;
wire nc18468;
wire nc18469;
wire nc18470;
wire nc18471;
wire nc18472;
wire nc18473;
wire nc18474;
wire nc18475;
wire nc18476;
wire nc18477;
wire nc18478;
wire nc18479;
wire nc18480;
wire nc18481;
wire nc18482;
wire nc18483;
wire nc18484;
wire nc18485;
wire nc18486;
wire nc18487;
wire nc18488;
wire nc18489;
wire nc18490;
wire nc18491;
wire nc18492;
wire nc18493;
wire nc18494;
wire nc18495;
wire nc18496;
wire nc18497;
wire nc18498;
wire nc18499;
wire nc18500;
wire nc18501;
wire nc18502;
wire nc18503;
wire nc18504;
wire nc18505;
wire nc18506;
wire nc18507;
wire nc18508;
wire nc18509;
wire nc18510;
wire nc18511;
wire nc18512;
wire nc18513;
wire nc18514;
wire nc18515;
wire nc18516;
wire nc18517;
wire nc18518;
wire nc18519;
wire nc18520;
wire nc18521;
wire nc18522;
wire nc18523;
wire nc18524;
wire nc18525;
wire nc18526;
wire nc18527;
wire nc18528;
wire nc18529;
wire nc18530;
wire nc18531;
wire nc18532;
wire nc18533;
wire nc18534;
wire nc18535;
wire nc18536;
wire nc18537;
wire nc18538;
wire nc18539;
wire nc18540;
wire nc18541;
wire nc18542;
wire nc18543;
wire nc18544;
wire nc18545;
wire nc18546;
wire nc18547;
wire nc18548;
wire nc18549;
wire nc18550;
wire nc18551;
wire nc18552;
wire nc18553;
wire nc18554;
wire nc18555;
wire nc18556;
wire nc18557;
wire nc18558;
wire nc18559;
wire nc18560;
wire nc18561;
wire nc18562;
wire nc18563;
wire nc18564;
wire nc18565;
wire nc18566;
wire nc18567;
wire nc18568;
wire nc18569;
wire nc18570;
wire nc18571;
wire nc18572;
wire nc18573;
wire nc18574;
wire nc18575;
wire nc18576;
wire nc18577;
wire nc18578;
wire nc18579;
wire nc18580;
wire nc18581;
wire nc18582;
wire nc18583;
wire nc18584;
wire nc18585;
wire nc18586;
wire nc18587;
wire nc18588;
wire nc18589;
wire nc18590;
wire nc18591;
wire nc18592;
wire nc18593;
wire nc18594;
wire nc18595;
wire nc18596;
wire nc18597;
wire nc18598;
wire nc18599;
wire nc18600;
wire nc18601;
wire nc18602;
wire nc18603;
wire nc18604;
wire nc18605;
wire nc18606;
wire nc18607;
wire nc18608;
wire nc18609;
wire nc18610;
wire nc18611;
wire nc18612;
wire nc18613;
wire nc18614;
wire nc18615;
wire nc18616;
wire nc18617;
wire nc18618;
wire nc18619;
wire nc18620;
wire nc18621;
wire nc18622;
wire nc18623;
wire nc18624;
wire nc18625;
wire nc18626;
wire nc18627;
wire nc18628;
wire nc18629;
wire nc18630;
wire nc18631;
wire nc18632;
wire nc18633;
wire nc18634;
wire nc18635;
wire nc18636;
wire nc18637;
wire nc18638;
wire nc18639;
wire nc18640;
wire nc18641;
wire nc18642;
wire nc18643;
wire nc18644;
wire nc18645;
wire nc18646;
wire nc18647;
wire nc18648;
wire nc18649;
wire nc18650;
wire nc18651;
wire nc18652;
wire nc18653;
wire nc18654;
wire nc18655;
wire nc18656;
wire nc18657;
wire nc18658;
wire nc18659;
wire nc18660;
wire nc18661;
wire nc18662;
wire nc18663;
wire nc18664;
wire nc18665;
wire nc18666;
wire nc18667;
wire nc18668;
wire nc18669;
wire nc18670;
wire nc18671;
wire nc18672;
wire nc18673;
wire nc18674;
wire nc18675;
wire nc18676;
wire nc18677;
wire nc18678;
wire nc18679;
wire nc18680;
wire nc18681;
wire nc18682;
wire nc18683;
wire nc18684;
wire nc18685;
wire nc18686;
wire nc18687;
wire nc18688;
wire nc18689;
wire nc18690;
wire nc18691;
wire nc18692;
wire nc18693;
wire nc18694;
wire nc18695;
wire nc18696;
wire nc18697;
wire nc18698;
wire nc18699;
wire nc18700;
wire nc18701;
wire nc18702;
wire nc18703;
wire nc18704;
wire nc18705;
wire nc18706;
wire nc18707;
wire nc18708;
wire nc18709;
wire nc18710;
wire nc18711;
wire nc18712;
wire nc18713;
wire nc18714;
wire nc18715;
wire nc18716;
wire nc18717;
wire nc18718;
wire nc18719;
wire nc18720;
wire nc18721;
wire nc18722;
wire nc18723;
wire nc18724;
wire nc18725;
wire nc18726;
wire nc18727;
wire nc18728;
wire nc18729;
wire nc18730;
wire nc18731;
wire nc18732;
wire nc18733;
wire nc18734;
wire nc18735;
wire nc18736;
wire nc18737;
wire nc18738;
wire nc18739;
wire nc18740;
wire nc18741;
wire nc18742;
wire nc18743;
wire nc18744;
wire nc18745;
wire nc18746;
wire nc18747;
wire nc18748;
wire nc18749;
wire nc18750;
wire nc18751;
wire nc18752;
wire nc18753;
wire nc18754;
wire nc18755;
wire nc18756;
wire nc18757;
wire nc18758;
wire nc18759;
wire nc18760;
wire nc18761;
wire nc18762;
wire nc18763;
wire nc18764;
wire nc18765;
wire nc18766;
wire nc18767;
wire nc18768;
wire nc18769;
wire nc18770;
wire nc18771;
wire nc18772;
wire nc18773;
wire nc18774;
wire nc18775;
wire nc18776;
wire nc18777;
wire nc18778;
wire nc18779;
wire nc18780;
wire nc18781;
wire nc18782;
wire nc18783;
wire nc18784;
wire nc18785;
wire nc18786;
wire nc18787;
wire nc18788;
wire nc18789;
wire nc18790;
wire nc18791;
wire nc18792;
wire nc18793;
wire nc18794;
wire nc18795;
wire nc18796;
wire nc18797;
wire nc18798;
wire nc18799;
wire nc18800;
wire nc18801;
wire nc18802;
wire nc18803;
wire nc18804;
wire nc18805;
wire nc18806;
wire nc18807;
wire nc18808;
wire nc18809;
wire nc18810;
wire nc18811;
wire nc18812;
wire nc18813;
wire nc18814;
wire nc18815;
wire nc18816;
wire nc18817;
wire nc18818;
wire nc18819;
wire nc18820;
wire nc18821;
wire nc18822;
wire nc18823;
wire nc18824;
wire nc18825;
wire nc18826;
wire nc18827;
wire nc18828;
wire nc18829;
wire nc18830;
wire nc18831;
wire nc18832;
wire nc18833;
wire nc18834;
wire nc18835;
wire nc18836;
wire nc18837;
wire nc18838;
wire nc18839;
wire nc18840;
wire nc18841;
wire nc18842;
wire nc18843;
wire nc18844;
wire nc18845;
wire nc18846;
wire nc18847;
wire nc18848;
wire nc18849;
wire nc18850;
wire nc18851;
wire nc18852;
wire nc18853;
wire nc18854;
wire nc18855;
wire nc18856;
wire nc18857;
wire nc18858;
wire nc18859;
wire nc18860;
wire nc18861;
wire nc18862;
wire nc18863;
wire nc18864;
wire nc18865;
wire nc18866;
wire nc18867;
wire nc18868;
wire nc18869;
wire nc18870;
wire nc18871;
wire nc18872;
wire nc18873;
wire nc18874;
wire nc18875;
wire nc18876;
wire nc18877;
wire nc18878;
wire nc18879;
wire nc18880;
wire nc18881;
wire nc18882;
wire nc18883;
wire nc18884;
wire nc18885;
wire nc18886;
wire nc18887;
wire nc18888;
wire nc18889;
wire nc18890;
wire nc18891;
wire nc18892;
wire nc18893;
wire nc18894;
wire nc18895;
wire nc18896;
wire nc18897;
wire nc18898;
wire nc18899;
wire nc18900;
wire nc18901;
wire nc18902;
wire nc18903;
wire nc18904;
wire nc18905;
wire nc18906;
wire nc18907;
wire nc18908;
wire nc18909;
wire nc18910;
wire nc18911;
wire nc18912;
wire nc18913;
wire nc18914;
wire nc18915;
wire nc18916;
wire nc18917;
wire nc18918;
wire nc18919;
wire nc18920;
wire nc18921;
wire nc18922;
wire nc18923;
wire nc18924;
wire nc18925;
wire nc18926;
wire nc18927;
wire nc18928;
wire nc18929;
wire nc18930;
wire nc18931;
wire nc18932;
wire nc18933;
wire nc18934;
wire nc18935;
wire nc18936;
wire nc18937;
wire nc18938;
wire nc18939;
wire nc18940;
wire nc18941;
wire nc18942;
wire nc18943;
wire nc18944;
wire nc18945;
wire nc18946;
wire nc18947;
wire nc18948;
wire nc18949;
wire nc18950;
wire nc18951;
wire nc18952;
wire nc18953;
wire nc18954;
wire nc18955;
wire nc18956;
wire nc18957;
wire nc18958;
wire nc18959;
wire nc18960;
wire nc18961;
wire nc18962;
wire nc18963;
wire nc18964;
wire nc18965;
wire nc18966;
wire nc18967;
wire nc18968;
wire nc18969;
wire nc18970;
wire nc18971;
wire nc18972;
wire nc18973;
wire nc18974;
wire nc18975;
wire nc18976;
wire nc18977;
wire nc18978;
wire nc18979;
wire nc18980;
wire nc18981;
wire nc18982;
wire nc18983;
wire nc18984;
wire nc18985;
wire nc18986;
wire nc18987;
wire nc18988;
wire nc18989;
wire nc18990;
wire nc18991;
wire nc18992;
wire nc18993;
wire nc18994;
wire nc18995;
wire nc18996;
wire nc18997;
wire nc18998;
wire nc18999;
wire nc19000;
wire nc19001;
wire nc19002;
wire nc19003;
wire nc19004;
wire nc19005;
wire nc19006;
wire nc19007;
wire nc19008;
wire nc19009;
wire nc19010;
wire nc19011;
wire nc19012;
wire nc19013;
wire nc19014;
wire nc19015;
wire nc19016;
wire nc19017;
wire nc19018;
wire nc19019;
wire nc19020;
wire nc19021;
wire nc19022;
wire nc19023;
wire nc19024;
wire nc19025;
wire nc19026;
wire nc19027;
wire nc19028;
wire nc19029;
wire nc19030;
wire nc19031;
wire nc19032;
wire nc19033;
wire nc19034;
wire nc19035;
wire nc19036;
wire nc19037;
wire nc19038;
wire nc19039;
wire nc19040;
wire nc19041;
wire nc19042;
wire nc19043;
wire nc19044;
wire nc19045;
wire nc19046;
wire nc19047;
wire nc19048;
wire nc19049;
wire nc19050;
wire nc19051;
wire nc19052;
wire nc19053;
wire nc19054;
wire nc19055;
wire nc19056;
wire nc19057;
wire nc19058;
wire nc19059;
wire nc19060;
wire nc19061;
wire nc19062;
wire nc19063;
wire nc19064;
wire nc19065;
wire nc19066;
wire nc19067;
wire nc19068;
wire nc19069;
wire nc19070;
wire nc19071;
wire nc19072;
wire nc19073;
wire nc19074;
wire nc19075;
wire nc19076;
wire nc19077;
wire nc19078;
wire nc19079;
wire nc19080;
wire nc19081;
wire nc19082;
wire nc19083;
wire nc19084;
wire nc19085;
wire nc19086;
wire nc19087;
wire nc19088;
wire nc19089;
wire nc19090;
wire nc19091;
wire nc19092;
wire nc19093;
wire nc19094;
wire nc19095;
wire nc19096;
wire nc19097;
wire nc19098;
wire nc19099;
wire nc19100;
wire nc19101;
wire nc19102;
wire nc19103;
wire nc19104;
wire nc19105;
wire nc19106;
wire nc19107;
wire nc19108;
wire nc19109;
wire nc19110;
wire nc19111;
wire nc19112;
wire nc19113;
wire nc19114;
wire nc19115;
wire nc19116;
wire nc19117;
wire nc19118;
wire nc19119;
wire nc19120;
wire nc19121;
wire nc19122;
wire nc19123;
wire nc19124;
wire nc19125;
wire nc19126;
wire nc19127;
wire nc19128;
wire nc19129;
wire nc19130;
wire nc19131;
wire nc19132;
wire nc19133;
wire nc19134;
wire nc19135;
wire nc19136;
wire nc19137;
wire nc19138;
wire nc19139;
wire nc19140;
wire nc19141;
wire nc19142;
wire nc19143;
wire nc19144;
wire nc19145;
wire nc19146;
wire nc19147;
wire nc19148;
wire nc19149;
wire nc19150;
wire nc19151;
wire nc19152;
wire nc19153;
wire nc19154;
wire nc19155;
wire nc19156;
wire nc19157;
wire nc19158;
wire nc19159;
wire nc19160;
wire nc19161;
wire nc19162;
wire nc19163;
wire nc19164;
wire nc19165;
wire nc19166;
wire nc19167;
wire nc19168;
wire nc19169;
wire nc19170;
wire nc19171;
wire nc19172;
wire nc19173;
wire nc19174;
wire nc19175;
wire nc19176;
wire nc19177;
wire nc19178;
wire nc19179;
wire nc19180;
wire nc19181;
wire nc19182;
wire nc19183;
wire nc19184;
wire nc19185;
wire nc19186;
wire nc19187;
wire nc19188;
wire nc19189;
wire nc19190;
wire nc19191;
wire nc19192;
wire nc19193;
wire nc19194;
wire nc19195;
wire nc19196;
wire nc19197;
wire nc19198;
wire nc19199;
wire nc19200;
wire nc19201;
wire nc19202;
wire nc19203;
wire nc19204;
wire nc19205;
wire nc19206;
wire nc19207;
wire nc19208;
wire nc19209;
wire nc19210;
wire nc19211;
wire nc19212;
wire nc19213;
wire nc19214;
wire nc19215;
wire nc19216;
wire nc19217;
wire nc19218;
wire nc19219;
wire nc19220;
wire nc19221;
wire nc19222;
wire nc19223;
wire nc19224;
wire nc19225;
wire nc19226;
wire nc19227;
wire nc19228;
wire nc19229;
wire nc19230;
wire nc19231;
wire nc19232;
wire nc19233;
wire nc19234;
wire nc19235;
wire nc19236;
wire nc19237;
wire nc19238;
wire nc19239;
wire nc19240;
wire nc19241;
wire nc19242;
wire nc19243;
wire nc19244;
wire nc19245;
wire nc19246;
wire nc19247;
wire nc19248;
wire nc19249;
wire nc19250;
wire nc19251;
wire nc19252;
wire nc19253;
wire nc19254;
wire nc19255;
wire nc19256;
wire nc19257;
wire nc19258;
wire nc19259;
wire nc19260;
wire nc19261;
wire nc19262;
wire nc19263;
wire nc19264;
wire nc19265;
wire nc19266;
wire nc19267;
wire nc19268;
wire nc19269;
wire nc19270;
wire nc19271;
wire nc19272;
wire nc19273;
wire nc19274;
wire nc19275;
wire nc19276;
wire nc19277;
wire nc19278;
wire nc19279;
wire nc19280;
wire nc19281;
wire nc19282;
wire nc19283;
wire nc19284;
wire nc19285;
wire nc19286;
wire nc19287;
wire nc19288;
wire nc19289;
wire nc19290;
wire nc19291;
wire nc19292;
wire nc19293;
wire nc19294;
wire nc19295;
wire nc19296;
wire nc19297;
wire nc19298;
wire nc19299;
wire nc19300;
wire nc19301;
wire nc19302;
wire nc19303;
wire nc19304;
wire nc19305;
wire nc19306;
wire nc19307;
wire nc19308;
wire nc19309;
wire nc19310;
wire nc19311;
wire nc19312;
wire nc19313;
wire nc19314;
wire nc19315;
wire nc19316;
wire nc19317;
wire nc19318;
wire nc19319;
wire nc19320;
wire nc19321;
wire nc19322;
wire nc19323;
wire nc19324;
wire nc19325;
wire nc19326;
wire nc19327;
wire nc19328;
wire nc19329;
wire nc19330;
wire nc19331;
wire nc19332;
wire nc19333;
wire nc19334;
wire nc19335;
wire nc19336;
wire nc19337;
wire nc19338;
wire nc19339;
wire nc19340;
wire nc19341;
wire nc19342;
wire nc19343;
wire nc19344;
wire nc19345;
wire nc19346;
wire nc19347;
wire nc19348;
wire nc19349;
wire nc19350;
wire nc19351;
wire nc19352;
wire nc19353;
wire nc19354;
wire nc19355;
wire nc19356;
wire nc19357;
wire nc19358;
wire nc19359;
wire nc19360;
wire nc19361;
wire nc19362;
wire nc19363;
wire nc19364;
wire nc19365;
wire nc19366;
wire nc19367;
wire nc19368;
wire nc19369;
wire nc19370;
wire nc19371;
wire nc19372;
wire nc19373;
wire nc19374;
wire nc19375;
wire nc19376;
wire nc19377;
wire nc19378;
wire nc19379;
wire nc19380;
wire nc19381;
wire nc19382;
wire nc19383;
wire nc19384;
wire nc19385;
wire nc19386;
wire nc19387;
wire nc19388;
wire nc19389;
wire nc19390;
wire nc19391;
wire nc19392;
wire nc19393;
wire nc19394;
wire nc19395;
wire nc19396;
wire nc19397;
wire nc19398;
wire nc19399;
wire nc19400;
wire nc19401;
wire nc19402;
wire nc19403;
wire nc19404;
wire nc19405;
wire nc19406;
wire nc19407;
wire nc19408;
wire nc19409;
wire nc19410;
wire nc19411;
wire nc19412;
wire nc19413;
wire nc19414;
wire nc19415;
wire nc19416;
wire nc19417;
wire nc19418;
wire nc19419;
wire nc19420;
wire nc19421;
wire nc19422;
wire nc19423;
wire nc19424;
wire nc19425;
wire nc19426;
wire nc19427;
wire nc19428;
wire nc19429;
wire nc19430;
wire nc19431;
wire nc19432;
wire nc19433;
wire nc19434;
wire nc19435;
wire nc19436;
wire nc19437;
wire nc19438;
wire nc19439;
wire nc19440;
wire nc19441;
wire nc19442;
wire nc19443;
wire nc19444;
wire nc19445;
wire nc19446;
wire nc19447;
wire nc19448;
wire nc19449;
wire nc19450;
wire nc19451;
wire nc19452;
wire nc19453;
wire nc19454;
wire nc19455;
wire nc19456;
wire nc19457;
wire nc19458;
wire nc19459;
wire nc19460;
wire nc19461;
wire nc19462;
wire nc19463;
wire nc19464;
wire nc19465;
wire nc19466;
wire nc19467;
wire nc19468;
wire nc19469;
wire nc19470;
wire nc19471;
wire nc19472;
wire nc19473;
wire nc19474;
wire nc19475;
wire nc19476;
wire nc19477;
wire nc19478;
wire nc19479;
wire nc19480;
wire nc19481;
wire nc19482;
wire nc19483;
wire nc19484;
wire nc19485;
wire nc19486;
wire nc19487;
wire nc19488;
wire nc19489;
wire nc19490;
wire nc19491;
wire nc19492;
wire nc19493;
wire nc19494;
wire nc19495;
wire nc19496;
wire nc19497;
wire nc19498;
wire nc19499;
wire nc19500;
wire nc19501;
wire nc19502;
wire nc19503;
wire nc19504;
wire nc19505;
wire nc19506;
wire nc19507;
wire nc19508;
wire nc19509;
wire nc19510;
wire nc19511;
wire nc19512;
wire nc19513;
wire nc19514;
wire nc19515;
wire nc19516;
wire nc19517;
wire nc19518;
wire nc19519;
wire nc19520;
wire nc19521;
wire nc19522;
wire nc19523;
wire nc19524;
wire nc19525;
wire nc19526;
wire nc19527;
wire nc19528;
wire nc19529;
wire nc19530;
wire nc19531;
wire nc19532;
wire nc19533;
wire nc19534;
wire nc19535;
wire nc19536;
wire nc19537;
wire nc19538;
wire nc19539;
wire nc19540;
wire nc19541;
wire nc19542;
wire nc19543;
wire nc19544;
wire nc19545;
wire nc19546;
wire nc19547;
wire nc19548;
wire nc19549;
wire nc19550;
wire nc19551;
wire nc19552;
wire nc19553;
wire nc19554;
wire nc19555;
wire nc19556;
wire nc19557;
wire nc19558;
wire nc19559;
wire nc19560;
wire nc19561;
wire nc19562;
wire nc19563;
wire nc19564;
wire nc19565;
wire nc19566;
wire nc19567;
wire nc19568;
wire nc19569;
wire nc19570;
wire nc19571;
wire nc19572;
wire nc19573;
wire nc19574;
wire nc19575;
wire nc19576;
wire nc19577;
wire nc19578;
wire nc19579;
wire nc19580;
wire nc19581;
wire nc19582;
wire nc19583;
wire nc19584;
wire nc19585;
wire nc19586;
wire nc19587;
wire nc19588;
wire nc19589;
wire nc19590;
wire nc19591;
wire nc19592;
wire nc19593;
wire nc19594;
wire nc19595;
wire nc19596;
wire nc19597;
wire nc19598;
wire nc19599;
wire nc19600;
wire nc19601;
wire nc19602;
wire nc19603;
wire nc19604;
wire nc19605;
wire nc19606;
wire nc19607;
wire nc19608;
wire nc19609;
wire nc19610;
wire nc19611;
wire nc19612;
wire nc19613;
wire nc19614;
wire nc19615;
wire nc19616;
wire nc19617;
wire nc19618;
wire nc19619;
wire nc19620;
wire nc19621;
wire nc19622;
wire nc19623;
wire nc19624;
wire nc19625;
wire nc19626;
wire nc19627;
wire nc19628;
wire nc19629;
wire nc19630;
wire nc19631;
wire nc19632;
wire nc19633;
wire nc19634;
wire nc19635;
wire nc19636;
wire nc19637;
wire nc19638;
wire nc19639;
wire nc19640;
wire nc19641;
wire nc19642;
wire nc19643;
wire nc19644;
wire nc19645;
wire nc19646;
wire nc19647;
wire nc19648;
wire nc19649;
wire nc19650;
wire nc19651;
wire nc19652;
wire nc19653;
wire nc19654;
wire nc19655;
wire nc19656;
wire nc19657;
wire nc19658;
wire nc19659;
wire nc19660;
wire nc19661;
wire nc19662;
wire nc19663;
wire nc19664;
wire nc19665;
wire nc19666;
wire nc19667;
wire nc19668;
wire nc19669;
wire nc19670;
wire nc19671;
wire nc19672;
wire nc19673;
wire nc19674;
wire nc19675;
wire nc19676;
wire nc19677;
wire nc19678;
wire nc19679;
wire nc19680;
wire nc19681;
wire nc19682;
wire nc19683;
wire nc19684;
wire nc19685;
wire nc19686;
wire nc19687;
wire nc19688;
wire nc19689;
wire nc19690;
wire nc19691;
wire nc19692;
wire nc19693;
wire nc19694;
wire nc19695;
wire nc19696;
wire nc19697;
wire nc19698;
wire nc19699;
wire nc19700;
wire nc19701;
wire nc19702;
wire nc19703;
wire nc19704;
wire nc19705;
wire nc19706;
wire nc19707;
wire nc19708;
wire nc19709;
wire nc19710;
wire nc19711;
wire nc19712;
wire nc19713;
wire nc19714;
wire nc19715;
wire nc19716;
wire nc19717;
wire nc19718;
wire nc19719;
wire nc19720;
wire nc19721;
wire nc19722;
wire nc19723;
wire nc19724;
wire nc19725;
wire nc19726;
wire nc19727;
wire nc19728;
wire nc19729;
wire nc19730;
wire nc19731;
wire nc19732;
wire nc19733;
wire nc19734;
wire nc19735;
wire nc19736;
wire nc19737;
wire nc19738;
wire nc19739;
wire nc19740;
wire nc19741;
wire nc19742;
wire nc19743;
wire nc19744;
wire nc19745;
wire nc19746;
wire nc19747;
wire nc19748;
wire nc19749;
wire nc19750;
wire nc19751;
wire nc19752;
wire nc19753;
wire nc19754;
wire nc19755;
wire nc19756;
wire nc19757;
wire nc19758;
wire nc19759;
wire nc19760;
wire nc19761;
wire nc19762;
wire nc19763;
wire nc19764;
wire nc19765;
wire nc19766;
wire nc19767;
wire nc19768;
wire nc19769;
wire nc19770;
wire nc19771;
wire nc19772;
wire nc19773;
wire nc19774;
wire nc19775;
wire nc19776;
wire nc19777;
wire nc19778;
wire nc19779;
wire nc19780;
wire nc19781;
wire nc19782;
wire nc19783;
wire nc19784;
wire nc19785;
wire nc19786;
wire nc19787;
wire nc19788;
wire nc19789;
wire nc19790;
wire nc19791;
wire nc19792;
wire nc19793;
wire nc19794;
wire nc19795;
wire nc19796;
wire nc19797;
wire nc19798;
wire nc19799;
wire nc19800;
wire nc19801;
wire nc19802;
wire nc19803;
wire nc19804;
wire nc19805;
wire nc19806;
wire nc19807;
wire nc19808;
wire nc19809;
wire nc19810;
wire nc19811;
wire nc19812;
wire nc19813;
wire nc19814;
wire nc19815;
wire nc19816;
wire nc19817;
wire nc19818;
wire nc19819;
wire nc19820;
wire nc19821;
wire nc19822;
wire nc19823;
wire nc19824;
wire nc19825;
wire nc19826;
wire nc19827;
wire nc19828;
wire nc19829;
wire nc19830;
wire nc19831;
wire nc19832;
wire nc19833;
wire nc19834;
wire nc19835;
wire nc19836;
wire nc19837;
wire nc19838;
wire nc19839;
wire nc19840;
wire nc19841;
wire nc19842;
wire nc19843;
wire nc19844;
wire nc19845;
wire nc19846;
wire nc19847;
wire nc19848;
wire nc19849;
wire nc19850;
wire nc19851;
wire nc19852;
wire nc19853;
wire nc19854;
wire nc19855;
wire nc19856;
wire nc19857;
wire nc19858;
wire nc19859;
wire nc19860;
wire nc19861;
wire nc19862;
wire nc19863;
wire nc19864;
wire nc19865;
wire nc19866;
wire nc19867;
wire nc19868;
wire nc19869;
wire nc19870;
wire nc19871;
wire nc19872;
wire nc19873;
wire nc19874;
wire nc19875;
wire nc19876;
wire nc19877;
wire nc19878;
wire nc19879;
wire nc19880;
wire nc19881;
wire nc19882;
wire nc19883;
wire nc19884;
wire nc19885;
wire nc19886;
wire nc19887;
wire nc19888;
wire nc19889;
wire nc19890;
wire nc19891;
wire nc19892;
wire nc19893;
wire nc19894;
wire nc19895;
wire nc19896;
wire nc19897;
wire nc19898;
wire nc19899;
wire nc19900;
wire nc19901;
wire nc19902;
wire nc19903;
wire nc19904;
wire nc19905;
wire nc19906;
wire nc19907;
wire nc19908;
wire nc19909;
wire nc19910;
wire nc19911;
wire nc19912;
wire nc19913;
wire nc19914;
wire nc19915;
wire nc19916;
wire nc19917;
wire nc19918;
wire nc19919;
wire nc19920;
wire nc19921;
wire nc19922;
wire nc19923;
wire nc19924;
wire nc19925;
wire nc19926;
wire nc19927;
wire nc19928;
wire nc19929;
wire nc19930;
wire nc19931;
wire nc19932;
wire nc19933;
wire nc19934;
wire nc19935;
wire nc19936;
wire nc19937;
wire nc19938;
wire nc19939;
wire nc19940;
wire nc19941;
wire nc19942;
wire nc19943;
wire nc19944;
wire nc19945;
wire nc19946;
wire nc19947;
wire nc19948;
wire nc19949;
wire nc19950;
wire nc19951;
wire nc19952;
wire nc19953;
wire nc19954;
wire nc19955;
wire nc19956;
wire nc19957;
wire nc19958;
wire nc19959;
wire nc19960;
wire nc19961;
wire nc19962;
wire nc19963;
wire nc19964;
wire nc19965;
wire nc19966;
wire nc19967;
wire nc19968;
wire nc19969;
wire nc19970;
wire nc19971;
wire nc19972;
wire nc19973;
wire nc19974;
wire nc19975;
wire nc19976;
wire nc19977;
wire nc19978;
wire nc19979;
wire nc19980;
wire nc19981;
wire nc19982;
wire nc19983;
wire nc19984;
wire nc19985;
wire nc19986;
wire nc19987;
wire nc19988;
wire nc19989;
wire nc19990;
wire nc19991;
wire nc19992;
wire nc19993;
wire nc19994;
wire nc19995;
wire nc19996;
wire nc19997;
wire nc19998;
wire nc19999;
wire nc20000;
wire nc20001;
wire nc20002;
wire nc20003;
wire nc20004;
wire nc20005;
wire nc20006;
wire nc20007;
wire nc20008;
wire nc20009;
wire nc20010;
wire nc20011;
wire nc20012;
wire nc20013;
wire nc20014;
wire nc20015;
wire nc20016;
wire nc20017;
wire nc20018;
wire nc20019;
wire nc20020;
wire nc20021;
wire nc20022;
wire nc20023;
wire nc20024;
wire nc20025;
wire nc20026;
wire nc20027;
wire nc20028;
wire nc20029;
wire nc20030;
wire nc20031;
wire nc20032;
wire nc20033;
wire nc20034;
wire nc20035;
wire nc20036;
wire nc20037;
wire nc20038;
wire nc20039;
wire nc20040;
wire nc20041;
wire nc20042;
wire nc20043;
wire nc20044;
wire nc20045;
wire nc20046;
wire nc20047;
wire nc20048;
wire nc20049;
wire nc20050;
wire nc20051;
wire nc20052;
wire nc20053;
wire nc20054;
wire nc20055;
wire nc20056;
wire nc20057;
wire nc20058;
wire nc20059;
wire nc20060;
wire nc20061;
wire nc20062;
wire nc20063;
wire nc20064;
wire nc20065;
wire nc20066;
wire nc20067;
wire nc20068;
wire nc20069;
wire nc20070;
wire nc20071;
wire nc20072;
wire nc20073;
wire nc20074;
wire nc20075;
wire nc20076;
wire nc20077;
wire nc20078;
wire nc20079;
wire nc20080;
wire nc20081;
wire nc20082;
wire nc20083;
wire nc20084;
wire nc20085;
wire nc20086;
wire nc20087;
wire nc20088;
wire nc20089;
wire nc20090;
wire nc20091;
wire nc20092;
wire nc20093;
wire nc20094;
wire nc20095;
wire nc20096;
wire nc20097;
wire nc20098;
wire nc20099;
wire nc20100;
wire nc20101;
wire nc20102;
wire nc20103;
wire nc20104;
wire nc20105;
wire nc20106;
wire nc20107;
wire nc20108;
wire nc20109;
wire nc20110;
wire nc20111;
wire nc20112;
wire nc20113;
wire nc20114;
wire nc20115;
wire nc20116;
wire nc20117;
wire nc20118;
wire nc20119;
wire nc20120;
wire nc20121;
wire nc20122;
wire nc20123;
wire nc20124;
wire nc20125;
wire nc20126;
wire nc20127;
wire nc20128;
wire nc20129;
wire nc20130;
wire nc20131;
wire nc20132;
wire nc20133;
wire nc20134;
wire nc20135;
wire nc20136;
wire nc20137;
wire nc20138;
wire nc20139;
wire nc20140;
wire nc20141;
wire nc20142;
wire nc20143;
wire nc20144;
wire nc20145;
wire nc20146;
wire nc20147;
wire nc20148;
wire nc20149;
wire nc20150;
wire nc20151;
wire nc20152;
wire nc20153;
wire nc20154;
wire nc20155;
wire nc20156;
wire nc20157;
wire nc20158;
wire nc20159;
wire nc20160;
wire nc20161;
wire nc20162;
wire nc20163;
wire nc20164;
wire nc20165;
wire nc20166;
wire nc20167;
wire nc20168;
wire nc20169;
wire nc20170;
wire nc20171;
wire nc20172;
wire nc20173;
wire nc20174;
wire nc20175;
wire nc20176;
wire nc20177;
wire nc20178;
wire nc20179;
wire nc20180;
wire nc20181;
wire nc20182;
wire nc20183;
wire nc20184;
wire nc20185;
wire nc20186;
wire nc20187;
wire nc20188;
wire nc20189;
wire nc20190;
wire nc20191;
wire nc20192;
wire nc20193;
wire nc20194;
wire nc20195;
wire nc20196;
wire nc20197;
wire nc20198;
wire nc20199;
wire nc20200;
wire nc20201;
wire nc20202;
wire nc20203;
wire nc20204;
wire nc20205;
wire nc20206;
wire nc20207;
wire nc20208;
wire nc20209;
wire nc20210;
wire nc20211;
wire nc20212;
wire nc20213;
wire nc20214;
wire nc20215;
wire nc20216;
wire nc20217;
wire nc20218;
wire nc20219;
wire nc20220;
wire nc20221;
wire nc20222;
wire nc20223;
wire nc20224;
wire nc20225;
wire nc20226;
wire nc20227;
wire nc20228;
wire nc20229;
wire nc20230;
wire nc20231;
wire nc20232;
wire nc20233;
wire nc20234;
wire nc20235;
wire nc20236;
wire nc20237;
wire nc20238;
wire nc20239;
wire nc20240;
wire nc20241;
wire nc20242;
wire nc20243;
wire nc20244;
wire nc20245;
wire nc20246;
wire nc20247;
wire nc20248;
wire nc20249;
wire nc20250;
wire nc20251;
wire nc20252;
wire nc20253;
wire nc20254;
wire nc20255;
wire nc20256;
wire nc20257;
wire nc20258;
wire nc20259;
wire nc20260;
wire nc20261;
wire nc20262;
wire nc20263;
wire nc20264;
wire nc20265;
wire nc20266;
wire nc20267;
wire nc20268;
wire nc20269;
wire nc20270;
wire nc20271;
wire nc20272;
wire nc20273;
wire nc20274;
wire nc20275;
wire nc20276;
wire nc20277;
wire nc20278;
wire nc20279;
wire nc20280;
wire nc20281;
wire nc20282;
wire nc20283;
wire nc20284;
wire nc20285;
wire nc20286;
wire nc20287;
wire nc20288;
wire nc20289;
wire nc20290;
wire nc20291;
wire nc20292;
wire nc20293;
wire nc20294;
wire nc20295;
wire nc20296;
wire nc20297;
wire nc20298;
wire nc20299;
wire nc20300;
wire nc20301;
wire nc20302;
wire nc20303;
wire nc20304;
wire nc20305;
wire nc20306;
wire nc20307;
wire nc20308;
wire nc20309;
wire nc20310;
wire nc20311;
wire nc20312;
wire nc20313;
wire nc20314;
wire nc20315;
wire nc20316;
wire nc20317;
wire nc20318;
wire nc20319;
wire nc20320;
wire nc20321;
wire nc20322;
wire nc20323;
wire nc20324;
wire nc20325;
wire nc20326;
wire nc20327;
wire nc20328;
wire nc20329;
wire nc20330;
wire nc20331;
wire nc20332;
wire nc20333;
wire nc20334;
wire nc20335;
wire nc20336;
wire nc20337;
wire nc20338;
wire nc20339;
wire nc20340;
wire nc20341;
wire nc20342;
wire nc20343;
wire nc20344;
wire nc20345;
wire nc20346;
wire nc20347;
wire nc20348;
wire nc20349;
wire nc20350;
wire nc20351;
wire nc20352;
wire nc20353;
wire nc20354;
wire nc20355;
wire nc20356;
wire nc20357;
wire nc20358;
wire nc20359;
wire nc20360;
wire nc20361;
wire nc20362;
wire nc20363;
wire nc20364;
wire nc20365;
wire nc20366;
wire nc20367;
wire nc20368;
wire nc20369;
wire nc20370;
wire nc20371;
wire nc20372;
wire nc20373;
wire nc20374;
wire nc20375;
wire nc20376;
wire nc20377;
wire nc20378;
wire nc20379;
wire nc20380;
wire nc20381;
wire nc20382;
wire nc20383;
wire nc20384;
wire nc20385;
wire nc20386;
wire nc20387;
wire nc20388;
wire nc20389;
wire nc20390;
wire nc20391;
wire nc20392;
wire nc20393;
wire nc20394;
wire nc20395;
wire nc20396;
wire nc20397;
wire nc20398;
wire nc20399;
wire nc20400;
wire nc20401;
wire nc20402;
wire nc20403;
wire nc20404;
wire nc20405;
wire nc20406;
wire nc20407;
wire nc20408;
wire nc20409;
wire nc20410;
wire nc20411;
wire nc20412;
wire nc20413;
wire nc20414;
wire nc20415;
wire nc20416;
wire nc20417;
wire nc20418;
wire nc20419;
wire nc20420;
wire nc20421;
wire nc20422;
wire nc20423;
wire nc20424;
wire nc20425;
wire nc20426;
wire nc20427;
wire nc20428;
wire nc20429;
wire nc20430;
wire nc20431;
wire nc20432;
wire nc20433;
wire nc20434;
wire nc20435;
wire nc20436;
wire nc20437;
wire nc20438;
wire nc20439;
wire nc20440;
wire nc20441;
wire nc20442;
wire nc20443;
wire nc20444;
wire nc20445;
wire nc20446;
wire nc20447;
wire nc20448;
wire nc20449;
wire nc20450;
wire nc20451;
wire nc20452;
wire nc20453;
wire nc20454;
wire nc20455;
wire nc20456;
wire nc20457;
wire nc20458;
wire nc20459;
wire nc20460;
wire nc20461;
wire nc20462;
wire nc20463;
wire nc20464;
wire nc20465;
wire nc20466;
wire nc20467;
wire nc20468;
wire nc20469;
wire nc20470;
wire nc20471;
wire nc20472;
wire nc20473;
wire nc20474;
wire nc20475;
wire nc20476;
wire nc20477;
wire nc20478;
wire nc20479;
wire nc20480;
wire nc20481;
wire nc20482;
wire nc20483;
wire nc20484;
wire nc20485;
wire nc20486;
wire nc20487;
wire nc20488;
wire nc20489;
wire nc20490;
wire nc20491;
wire nc20492;
wire nc20493;
wire nc20494;
wire nc20495;
wire nc20496;
wire nc20497;
wire nc20498;
wire nc20499;
wire nc20500;
wire nc20501;
wire nc20502;
wire nc20503;
wire nc20504;
wire nc20505;
wire nc20506;
wire nc20507;
wire nc20508;
wire nc20509;
wire nc20510;
wire nc20511;
wire nc20512;
wire nc20513;
wire nc20514;
wire nc20515;
wire nc20516;
wire nc20517;
wire nc20518;
wire nc20519;
wire nc20520;
wire nc20521;
wire nc20522;
wire nc20523;
wire nc20524;
wire nc20525;
wire nc20526;
wire nc20527;
wire nc20528;
wire nc20529;
wire nc20530;
wire nc20531;
wire nc20532;
wire nc20533;
wire nc20534;
wire nc20535;
wire nc20536;
wire nc20537;
wire nc20538;
wire nc20539;
wire nc20540;
wire nc20541;
wire nc20542;
wire nc20543;
wire nc20544;
wire nc20545;
wire nc20546;
wire nc20547;
wire nc20548;
wire nc20549;
wire nc20550;
wire nc20551;
wire nc20552;
wire nc20553;
wire nc20554;
wire nc20555;
wire nc20556;
wire nc20557;
wire nc20558;
wire nc20559;
wire nc20560;
wire nc20561;
wire nc20562;
wire nc20563;
wire nc20564;
wire nc20565;
wire nc20566;
wire nc20567;
wire nc20568;
wire nc20569;
wire nc20570;
wire nc20571;
wire nc20572;
wire nc20573;
wire nc20574;
wire nc20575;
wire nc20576;
wire nc20577;
wire nc20578;
wire nc20579;
wire nc20580;
wire nc20581;
wire nc20582;
wire nc20583;
wire nc20584;
wire nc20585;
wire nc20586;
wire nc20587;
wire nc20588;
wire nc20589;
wire nc20590;
wire nc20591;
wire nc20592;
wire nc20593;
wire nc20594;
wire nc20595;
wire nc20596;
wire nc20597;
wire nc20598;
wire nc20599;
wire nc20600;
wire nc20601;
wire nc20602;
wire nc20603;
wire nc20604;
wire nc20605;
wire nc20606;
wire nc20607;
wire nc20608;
wire nc20609;
wire nc20610;
wire nc20611;
wire nc20612;
wire nc20613;
wire nc20614;
wire nc20615;
wire nc20616;
wire nc20617;
wire nc20618;
wire nc20619;
wire nc20620;
wire nc20621;
wire nc20622;
wire nc20623;
wire nc20624;
wire nc20625;
wire nc20626;
wire nc20627;
wire nc20628;
wire nc20629;
wire nc20630;
wire nc20631;
wire nc20632;
wire nc20633;
wire nc20634;
wire nc20635;
wire nc20636;
wire nc20637;
wire nc20638;
wire nc20639;
wire nc20640;
wire nc20641;
wire nc20642;
wire nc20643;
wire nc20644;
wire nc20645;
wire nc20646;
wire nc20647;
wire nc20648;
wire nc20649;
wire nc20650;
wire nc20651;
wire nc20652;
wire nc20653;
wire nc20654;
wire nc20655;
wire nc20656;
wire nc20657;
wire nc20658;
wire nc20659;
wire nc20660;
wire nc20661;
wire nc20662;
wire nc20663;
wire nc20664;
wire nc20665;
wire nc20666;
wire nc20667;
wire nc20668;
wire nc20669;
wire nc20670;
wire nc20671;
wire nc20672;
wire nc20673;
wire nc20674;
wire nc20675;
wire nc20676;
wire nc20677;
wire nc20678;
wire nc20679;
wire nc20680;
wire nc20681;
wire nc20682;
wire nc20683;
wire nc20684;
wire nc20685;
wire nc20686;
wire nc20687;
wire nc20688;
wire nc20689;
wire nc20690;
wire nc20691;
wire nc20692;
wire nc20693;
wire nc20694;
wire nc20695;
wire nc20696;
wire nc20697;
wire nc20698;
wire nc20699;
wire nc20700;
wire nc20701;
wire nc20702;
wire nc20703;
wire nc20704;
wire nc20705;
wire nc20706;
wire nc20707;
wire nc20708;
wire nc20709;
wire nc20710;
wire nc20711;
wire nc20712;
wire nc20713;
wire nc20714;
wire nc20715;
wire nc20716;
wire nc20717;
wire nc20718;
wire nc20719;
wire nc20720;
wire nc20721;
wire nc20722;
wire nc20723;
wire nc20724;
wire nc20725;
wire nc20726;
wire nc20727;
wire nc20728;
wire nc20729;
wire nc20730;
wire nc20731;
wire nc20732;
wire nc20733;
wire nc20734;
wire nc20735;
wire nc20736;
wire nc20737;
wire nc20738;
wire nc20739;
wire nc20740;
wire nc20741;
wire nc20742;
wire nc20743;
wire nc20744;
wire nc20745;
wire nc20746;
wire nc20747;
wire nc20748;
wire nc20749;
wire nc20750;
wire nc20751;
wire nc20752;
wire nc20753;
wire nc20754;
wire nc20755;
wire nc20756;
wire nc20757;
wire nc20758;
wire nc20759;
wire nc20760;
wire nc20761;
wire nc20762;
wire nc20763;
wire nc20764;
wire nc20765;
wire nc20766;
wire nc20767;
wire nc20768;
wire nc20769;
wire nc20770;
wire nc20771;
wire nc20772;
wire nc20773;
wire nc20774;
wire nc20775;
wire nc20776;
wire nc20777;
wire nc20778;
wire nc20779;
wire nc20780;
wire nc20781;
wire nc20782;
wire nc20783;
wire nc20784;
wire nc20785;
wire nc20786;
wire nc20787;
wire nc20788;
wire nc20789;
wire nc20790;
wire nc20791;
wire nc20792;
wire nc20793;
wire nc20794;
wire nc20795;
wire nc20796;
wire nc20797;
wire nc20798;
wire nc20799;
wire nc20800;
wire nc20801;
wire nc20802;
wire nc20803;
wire nc20804;
wire nc20805;
wire nc20806;
wire nc20807;
wire nc20808;
wire nc20809;
wire nc20810;
wire nc20811;
wire nc20812;
wire nc20813;
wire nc20814;
wire nc20815;
wire nc20816;
wire nc20817;
wire nc20818;
wire nc20819;
wire nc20820;
wire nc20821;
wire nc20822;
wire nc20823;
wire nc20824;
wire nc20825;
wire nc20826;
wire nc20827;
wire nc20828;
wire nc20829;
wire nc20830;
wire nc20831;
wire nc20832;
wire nc20833;
wire nc20834;
wire nc20835;
wire nc20836;
wire nc20837;
wire nc20838;
wire nc20839;
wire nc20840;
wire nc20841;
wire nc20842;
wire nc20843;
wire nc20844;
wire nc20845;
wire nc20846;
wire nc20847;
wire nc20848;
wire nc20849;
wire nc20850;
wire nc20851;
wire nc20852;
wire nc20853;
wire nc20854;
wire nc20855;
wire nc20856;
wire nc20857;
wire nc20858;
wire nc20859;
wire nc20860;
wire nc20861;
wire nc20862;
wire nc20863;
wire nc20864;
wire nc20865;
wire nc20866;
wire nc20867;
wire nc20868;
wire nc20869;
wire nc20870;
wire nc20871;
wire nc20872;
wire nc20873;
wire nc20874;
wire nc20875;
wire nc20876;
wire nc20877;
wire nc20878;
wire nc20879;
wire nc20880;
wire nc20881;
wire nc20882;
wire nc20883;
wire nc20884;
wire nc20885;
wire nc20886;
wire nc20887;
wire nc20888;
wire nc20889;
wire nc20890;
wire nc20891;
wire nc20892;
wire nc20893;
wire nc20894;
wire nc20895;
wire nc20896;
wire nc20897;
wire nc20898;
wire nc20899;
wire nc20900;
wire nc20901;
wire nc20902;
wire nc20903;
wire nc20904;
wire nc20905;
wire nc20906;
wire nc20907;
wire nc20908;
wire nc20909;
wire nc20910;
wire nc20911;
wire nc20912;
wire nc20913;
wire nc20914;
wire nc20915;
wire nc20916;
wire nc20917;
wire nc20918;
wire nc20919;
wire nc20920;
wire nc20921;
wire nc20922;
wire nc20923;
wire nc20924;
wire nc20925;
wire nc20926;
wire nc20927;
wire nc20928;
wire nc20929;
wire nc20930;
wire nc20931;
wire nc20932;
wire nc20933;
wire nc20934;
wire nc20935;
wire nc20936;
wire nc20937;
wire nc20938;
wire nc20939;
wire nc20940;
wire nc20941;
wire nc20942;
wire nc20943;
wire nc20944;
wire nc20945;
wire nc20946;
wire nc20947;
wire nc20948;
wire nc20949;
wire nc20950;
wire nc20951;
wire nc20952;
wire nc20953;
wire nc20954;
wire nc20955;
wire nc20956;
wire nc20957;
wire nc20958;
wire nc20959;
wire nc20960;
wire nc20961;
wire nc20962;
wire nc20963;
wire nc20964;
wire nc20965;
wire nc20966;
wire nc20967;
wire nc20968;
wire nc20969;
wire nc20970;
wire nc20971;
wire nc20972;
wire nc20973;
wire nc20974;
wire nc20975;
wire nc20976;
wire nc20977;
wire nc20978;
wire nc20979;
wire nc20980;
wire nc20981;
wire nc20982;
wire nc20983;
wire nc20984;
wire nc20985;
wire nc20986;
wire nc20987;
wire nc20988;
wire nc20989;
wire nc20990;
wire nc20991;
wire nc20992;
wire nc20993;
wire nc20994;
wire nc20995;
wire nc20996;
wire nc20997;
wire nc20998;
wire nc20999;
wire nc21000;
wire nc21001;
wire nc21002;
wire nc21003;
wire nc21004;
wire nc21005;
wire nc21006;
wire nc21007;
wire nc21008;
wire nc21009;
wire nc21010;
wire nc21011;
wire nc21012;
wire nc21013;
wire nc21014;
wire nc21015;
wire nc21016;
wire nc21017;
wire nc21018;
wire nc21019;
wire nc21020;
wire nc21021;
wire nc21022;
wire nc21023;
wire nc21024;
wire nc21025;
wire nc21026;
wire nc21027;
wire nc21028;
wire nc21029;
wire nc21030;
wire nc21031;
wire nc21032;
wire nc21033;
wire nc21034;
wire nc21035;
wire nc21036;
wire nc21037;
wire nc21038;
wire nc21039;
wire nc21040;
wire nc21041;
wire nc21042;
wire nc21043;
wire nc21044;
wire nc21045;
wire nc21046;
wire nc21047;
wire nc21048;
wire nc21049;
wire nc21050;
wire nc21051;
wire nc21052;
wire nc21053;
wire nc21054;
wire nc21055;
wire nc21056;
wire nc21057;
wire nc21058;
wire nc21059;
wire nc21060;
wire nc21061;
wire nc21062;
wire nc21063;
wire nc21064;
wire nc21065;
wire nc21066;
wire nc21067;
wire nc21068;
wire nc21069;
wire nc21070;
wire nc21071;
wire nc21072;
wire nc21073;
wire nc21074;
wire nc21075;
wire nc21076;
wire nc21077;
wire nc21078;
wire nc21079;
wire nc21080;
wire nc21081;
wire nc21082;
wire nc21083;
wire nc21084;
wire nc21085;
wire nc21086;
wire nc21087;
wire nc21088;
wire nc21089;
wire nc21090;
wire nc21091;
wire nc21092;
wire nc21093;
wire nc21094;
wire nc21095;
wire nc21096;
wire nc21097;
wire nc21098;
wire nc21099;
wire nc21100;
wire nc21101;
wire nc21102;
wire nc21103;
wire nc21104;
wire nc21105;
wire nc21106;
wire nc21107;
wire nc21108;
wire nc21109;
wire nc21110;
wire nc21111;
wire nc21112;
wire nc21113;
wire nc21114;
wire nc21115;
wire nc21116;
wire nc21117;
wire nc21118;
wire nc21119;
wire nc21120;
wire nc21121;
wire nc21122;
wire nc21123;
wire nc21124;
wire nc21125;
wire nc21126;
wire nc21127;
wire nc21128;
wire nc21129;
wire nc21130;
wire nc21131;
wire nc21132;
wire nc21133;
wire nc21134;
wire nc21135;
wire nc21136;
wire nc21137;
wire nc21138;
wire nc21139;
wire nc21140;
wire nc21141;
wire nc21142;
wire nc21143;
wire nc21144;
wire nc21145;
wire nc21146;
wire nc21147;
wire nc21148;
wire nc21149;
wire nc21150;
wire nc21151;
wire nc21152;
wire nc21153;
wire nc21154;
wire nc21155;
wire nc21156;
wire nc21157;
wire nc21158;
wire nc21159;
wire nc21160;
wire nc21161;
wire nc21162;
wire nc21163;
wire nc21164;
wire nc21165;
wire nc21166;
wire nc21167;
wire nc21168;
wire nc21169;
wire nc21170;
wire nc21171;
wire nc21172;
wire nc21173;
wire nc21174;
wire nc21175;
wire nc21176;
wire nc21177;
wire nc21178;
wire nc21179;
wire nc21180;
wire nc21181;
wire nc21182;
wire nc21183;
wire nc21184;
wire nc21185;
wire nc21186;
wire nc21187;
wire nc21188;
wire nc21189;
wire nc21190;
wire nc21191;
wire nc21192;
wire nc21193;
wire nc21194;
wire nc21195;
wire nc21196;
wire nc21197;
wire nc21198;
wire nc21199;
wire nc21200;
wire nc21201;
wire nc21202;
wire nc21203;
wire nc21204;
wire nc21205;
wire nc21206;
wire nc21207;
wire nc21208;
wire nc21209;
wire nc21210;
wire nc21211;
wire nc21212;
wire nc21213;
wire nc21214;
wire nc21215;
wire nc21216;
wire nc21217;
wire nc21218;
wire nc21219;
wire nc21220;
wire nc21221;
wire nc21222;
wire nc21223;
wire nc21224;
wire nc21225;
wire nc21226;
wire nc21227;
wire nc21228;
wire nc21229;
wire nc21230;
wire nc21231;
wire nc21232;
wire nc21233;
wire nc21234;
wire nc21235;
wire nc21236;
wire nc21237;
wire nc21238;
wire nc21239;
wire nc21240;
wire nc21241;
wire nc21242;
wire nc21243;
wire nc21244;
wire nc21245;
wire nc21246;
wire nc21247;
wire nc21248;
wire nc21249;
wire nc21250;
wire nc21251;
wire nc21252;
wire nc21253;
wire nc21254;
wire nc21255;
wire nc21256;
wire nc21257;
wire nc21258;
wire nc21259;
wire nc21260;
wire nc21261;
wire nc21262;
wire nc21263;
wire nc21264;
wire nc21265;
wire nc21266;
wire nc21267;
wire nc21268;
wire nc21269;
wire nc21270;
wire nc21271;
wire nc21272;
wire nc21273;
wire nc21274;
wire nc21275;
wire nc21276;
wire nc21277;
wire nc21278;
wire nc21279;
wire nc21280;
wire nc21281;
wire nc21282;
wire nc21283;
wire nc21284;
wire nc21285;
wire nc21286;
wire nc21287;
wire nc21288;
wire nc21289;
wire nc21290;
wire nc21291;
wire nc21292;
wire nc21293;
wire nc21294;
wire nc21295;
wire nc21296;
wire nc21297;
wire nc21298;
wire nc21299;
wire nc21300;
wire nc21301;
wire nc21302;
wire nc21303;
wire nc21304;
wire nc21305;
wire nc21306;
wire nc21307;
wire nc21308;
wire nc21309;
wire nc21310;
wire nc21311;
wire nc21312;
wire nc21313;
wire nc21314;
wire nc21315;
wire nc21316;
wire nc21317;
wire nc21318;
wire nc21319;
wire nc21320;
wire nc21321;
wire nc21322;
wire nc21323;
wire nc21324;
wire nc21325;
wire nc21326;
wire nc21327;
wire nc21328;
wire nc21329;
wire nc21330;
wire nc21331;
wire nc21332;
wire nc21333;
wire nc21334;
wire nc21335;
wire nc21336;
wire nc21337;
wire nc21338;
wire nc21339;
wire nc21340;
wire nc21341;
wire nc21342;
wire nc21343;
wire nc21344;
wire nc21345;
wire nc21346;
wire nc21347;
wire nc21348;
wire nc21349;
wire nc21350;
wire nc21351;
wire nc21352;
wire nc21353;
wire nc21354;
wire nc21355;
wire nc21356;
wire nc21357;
wire nc21358;
wire nc21359;
wire nc21360;
wire nc21361;
wire nc21362;
wire nc21363;
wire nc21364;
wire nc21365;
wire nc21366;
wire nc21367;
wire nc21368;
wire nc21369;
wire nc21370;
wire nc21371;
wire nc21372;
wire nc21373;
wire nc21374;
wire nc21375;
wire nc21376;
wire nc21377;
wire nc21378;
wire nc21379;
wire nc21380;
wire nc21381;
wire nc21382;
wire nc21383;
wire nc21384;
wire nc21385;
wire nc21386;
wire nc21387;
wire nc21388;
wire nc21389;
wire nc21390;
wire nc21391;
wire nc21392;
wire nc21393;
wire nc21394;
wire nc21395;
wire nc21396;
wire nc21397;
wire nc21398;
wire nc21399;
wire nc21400;
wire nc21401;
wire nc21402;
wire nc21403;
wire nc21404;
wire nc21405;
wire nc21406;
wire nc21407;
wire nc21408;
wire nc21409;
wire nc21410;
wire nc21411;
wire nc21412;
wire nc21413;
wire nc21414;
wire nc21415;
wire nc21416;
wire nc21417;
wire nc21418;
wire nc21419;
wire nc21420;
wire nc21421;
wire nc21422;
wire nc21423;
wire nc21424;
wire nc21425;
wire nc21426;
wire nc21427;
wire nc21428;
wire nc21429;
wire nc21430;
wire nc21431;
wire nc21432;
wire nc21433;
wire nc21434;
wire nc21435;
wire nc21436;
wire nc21437;
wire nc21438;
wire nc21439;
wire nc21440;
wire nc21441;
wire nc21442;
wire nc21443;
wire nc21444;
wire nc21445;
wire nc21446;
wire nc21447;
wire nc21448;
wire nc21449;
wire nc21450;
wire nc21451;
wire nc21452;
wire nc21453;
wire nc21454;
wire nc21455;
wire nc21456;
wire nc21457;
wire nc21458;
wire nc21459;
wire nc21460;
wire nc21461;
wire nc21462;
wire nc21463;
wire nc21464;
wire nc21465;
wire nc21466;
wire nc21467;
wire nc21468;
wire nc21469;
wire nc21470;
wire nc21471;
wire nc21472;
wire nc21473;
wire nc21474;
wire nc21475;
wire nc21476;
wire nc21477;
wire nc21478;
wire nc21479;
wire nc21480;
wire nc21481;
wire nc21482;
wire nc21483;
wire nc21484;
wire nc21485;
wire nc21486;
wire nc21487;
wire nc21488;
wire nc21489;
wire nc21490;
wire nc21491;
wire nc21492;
wire nc21493;
wire nc21494;
wire nc21495;
wire nc21496;
wire nc21497;
wire nc21498;
wire nc21499;
wire nc21500;
wire nc21501;
wire nc21502;
wire nc21503;
wire nc21504;
wire nc21505;
wire nc21506;
wire nc21507;
wire nc21508;
wire nc21509;
wire nc21510;
wire nc21511;
wire nc21512;
wire nc21513;
wire nc21514;
wire nc21515;
wire nc21516;
wire nc21517;
wire nc21518;
wire nc21519;
wire nc21520;
wire nc21521;
wire nc21522;
wire nc21523;
wire nc21524;
wire nc21525;
wire nc21526;
wire nc21527;
wire nc21528;
wire nc21529;
wire nc21530;
wire nc21531;
wire nc21532;
wire nc21533;
wire nc21534;
wire nc21535;
wire nc21536;
wire nc21537;
wire nc21538;
wire nc21539;
wire nc21540;
wire nc21541;
wire nc21542;
wire nc21543;
wire nc21544;
wire nc21545;
wire nc21546;
wire nc21547;
wire nc21548;
wire nc21549;
wire nc21550;
wire nc21551;
wire nc21552;
wire nc21553;
wire nc21554;
wire nc21555;
wire nc21556;
wire nc21557;
wire nc21558;
wire nc21559;
wire nc21560;
wire nc21561;
wire nc21562;
wire nc21563;
wire nc21564;
wire nc21565;
wire nc21566;
wire nc21567;
wire nc21568;
wire nc21569;
wire nc21570;
wire nc21571;
wire nc21572;
wire nc21573;
wire nc21574;
wire nc21575;
wire nc21576;
wire nc21577;
wire nc21578;
wire nc21579;
wire nc21580;
wire nc21581;
wire nc21582;
wire nc21583;
wire nc21584;
wire nc21585;
wire nc21586;
wire nc21587;
wire nc21588;
wire nc21589;
wire nc21590;
wire nc21591;
wire nc21592;
wire nc21593;
wire nc21594;
wire nc21595;
wire nc21596;
wire nc21597;
wire nc21598;
wire nc21599;
wire nc21600;
wire nc21601;
wire nc21602;
wire nc21603;
wire nc21604;
wire nc21605;
wire nc21606;
wire nc21607;
wire nc21608;
wire nc21609;
wire nc21610;
wire nc21611;
wire nc21612;
wire nc21613;
wire nc21614;
wire nc21615;
wire nc21616;
wire nc21617;
wire nc21618;
wire nc21619;
wire nc21620;
wire nc21621;
wire nc21622;
wire nc21623;
wire nc21624;
wire nc21625;
wire nc21626;
wire nc21627;
wire nc21628;
wire nc21629;
wire nc21630;
wire nc21631;
wire nc21632;
wire nc21633;
wire nc21634;
wire nc21635;
wire nc21636;
wire nc21637;
wire nc21638;
wire nc21639;
wire nc21640;
wire nc21641;
wire nc21642;
wire nc21643;
wire nc21644;
wire nc21645;
wire nc21646;
wire nc21647;
wire nc21648;
wire nc21649;
wire nc21650;
wire nc21651;
wire nc21652;
wire nc21653;
wire nc21654;
wire nc21655;
wire nc21656;
wire nc21657;
wire nc21658;
wire nc21659;
wire nc21660;
wire nc21661;
wire nc21662;
wire nc21663;
wire nc21664;
wire nc21665;
wire nc21666;
wire nc21667;
wire nc21668;
wire nc21669;
wire nc21670;
wire nc21671;
wire nc21672;
wire nc21673;
wire nc21674;
wire nc21675;
wire nc21676;
wire nc21677;
wire nc21678;
wire nc21679;
wire nc21680;
wire nc21681;
wire nc21682;
wire nc21683;
wire nc21684;
wire nc21685;
wire nc21686;
wire nc21687;
wire nc21688;
wire nc21689;
wire nc21690;
wire nc21691;
wire nc21692;
wire nc21693;
wire nc21694;
wire nc21695;
wire nc21696;
wire nc21697;
wire nc21698;
wire nc21699;
wire nc21700;
wire nc21701;
wire nc21702;
wire nc21703;
wire nc21704;
wire nc21705;
wire nc21706;
wire nc21707;
wire nc21708;
wire nc21709;
wire nc21710;
wire nc21711;
wire nc21712;
wire nc21713;
wire nc21714;
wire nc21715;
wire nc21716;
wire nc21717;
wire nc21718;
wire nc21719;
wire nc21720;
wire nc21721;
wire nc21722;
wire nc21723;
wire nc21724;
wire nc21725;
wire nc21726;
wire nc21727;
wire nc21728;
wire nc21729;
wire nc21730;
wire nc21731;
wire nc21732;
wire nc21733;
wire nc21734;
wire nc21735;
wire nc21736;
wire nc21737;
wire nc21738;
wire nc21739;
wire nc21740;
wire nc21741;
wire nc21742;
wire nc21743;
wire nc21744;
wire nc21745;
wire nc21746;
wire nc21747;
wire nc21748;
wire nc21749;
wire nc21750;
wire nc21751;
wire nc21752;
wire nc21753;
wire nc21754;
wire nc21755;
wire nc21756;
wire nc21757;
wire nc21758;
wire nc21759;
wire nc21760;
wire nc21761;
wire nc21762;
wire nc21763;
wire nc21764;
wire nc21765;
wire nc21766;
wire nc21767;
wire nc21768;
wire nc21769;
wire nc21770;
wire nc21771;
wire nc21772;
wire nc21773;
wire nc21774;
wire nc21775;
wire nc21776;
wire nc21777;
wire nc21778;
wire nc21779;
wire nc21780;
wire nc21781;
wire nc21782;
wire nc21783;
wire nc21784;
wire nc21785;
wire nc21786;
wire nc21787;
wire nc21788;
wire nc21789;
wire nc21790;
wire nc21791;
wire nc21792;
wire nc21793;
wire nc21794;
wire nc21795;
wire nc21796;
wire nc21797;
wire nc21798;
wire nc21799;
wire nc21800;
wire nc21801;
wire nc21802;
wire nc21803;
wire nc21804;
wire nc21805;
wire nc21806;
wire nc21807;
wire nc21808;
wire nc21809;
wire nc21810;
wire nc21811;
wire nc21812;
wire nc21813;
wire nc21814;
wire nc21815;
wire nc21816;
wire nc21817;
wire nc21818;
wire nc21819;
wire nc21820;
wire nc21821;
wire nc21822;
wire nc21823;
wire nc21824;
wire nc21825;
wire nc21826;
wire nc21827;
wire nc21828;
wire nc21829;
wire nc21830;
wire nc21831;
wire nc21832;
wire nc21833;
wire nc21834;
wire nc21835;
wire nc21836;
wire nc21837;
wire nc21838;
wire nc21839;
wire nc21840;
wire nc21841;
wire nc21842;
wire nc21843;
wire nc21844;
wire nc21845;
wire nc21846;
wire nc21847;
wire nc21848;
wire nc21849;
wire nc21850;
wire nc21851;
wire nc21852;
wire nc21853;
wire nc21854;
wire nc21855;
wire nc21856;
wire nc21857;
wire nc21858;
wire nc21859;
wire nc21860;
wire nc21861;
wire nc21862;
wire nc21863;
wire nc21864;
wire nc21865;
wire nc21866;
wire nc21867;
wire nc21868;
wire nc21869;
wire nc21870;
wire nc21871;
wire nc21872;
wire nc21873;
wire nc21874;
wire nc21875;
wire nc21876;
wire nc21877;
wire nc21878;
wire nc21879;
wire nc21880;
wire nc21881;
wire nc21882;
wire nc21883;
wire nc21884;
wire nc21885;
wire nc21886;
wire nc21887;
wire nc21888;
wire nc21889;
wire nc21890;
wire nc21891;
wire nc21892;
wire nc21893;
wire nc21894;
wire nc21895;
wire nc21896;
wire nc21897;
wire nc21898;
wire nc21899;
wire nc21900;
wire nc21901;
wire nc21902;
wire nc21903;
wire nc21904;
wire nc21905;
wire nc21906;
wire nc21907;
wire nc21908;
wire nc21909;
wire nc21910;
wire nc21911;
wire nc21912;
wire nc21913;
wire nc21914;
wire nc21915;
wire nc21916;
wire nc21917;
wire nc21918;
wire nc21919;
wire nc21920;
wire nc21921;
wire nc21922;
wire nc21923;
wire nc21924;
wire nc21925;
wire nc21926;
wire nc21927;
wire nc21928;
wire nc21929;
wire nc21930;
wire nc21931;
wire nc21932;
wire nc21933;
wire nc21934;
wire nc21935;
wire nc21936;
wire nc21937;
wire nc21938;
wire nc21939;
wire nc21940;
wire nc21941;
wire nc21942;
wire nc21943;
wire nc21944;
wire nc21945;
wire nc21946;
wire nc21947;
wire nc21948;
wire nc21949;
wire nc21950;
wire nc21951;
wire nc21952;
wire nc21953;
wire nc21954;
wire nc21955;
wire nc21956;
wire nc21957;
wire nc21958;
wire nc21959;
wire nc21960;
wire nc21961;
wire nc21962;
wire nc21963;
wire nc21964;
wire nc21965;
wire nc21966;
wire nc21967;
wire nc21968;
wire nc21969;
wire nc21970;
wire nc21971;
wire nc21972;
wire nc21973;
wire nc21974;
wire nc21975;
wire nc21976;
wire nc21977;
wire nc21978;
wire nc21979;
wire nc21980;
wire nc21981;
wire nc21982;
wire nc21983;
wire nc21984;
wire nc21985;
wire nc21986;
wire nc21987;
wire nc21988;
wire nc21989;
wire nc21990;
wire nc21991;
wire nc21992;
wire nc21993;
wire nc21994;
wire nc21995;
wire nc21996;
wire nc21997;
wire nc21998;
wire nc21999;
wire nc22000;
wire nc22001;
wire nc22002;
wire nc22003;
wire nc22004;
wire nc22005;
wire nc22006;
wire nc22007;
wire nc22008;
wire nc22009;
wire nc22010;
wire nc22011;
wire nc22012;
wire nc22013;
wire nc22014;
wire nc22015;
wire nc22016;
wire nc22017;
wire nc22018;
wire nc22019;
wire nc22020;
wire nc22021;
wire nc22022;
wire nc22023;
wire nc22024;
wire nc22025;
wire nc22026;
wire nc22027;
wire nc22028;
wire nc22029;
wire nc22030;
wire nc22031;
wire nc22032;
wire nc22033;
wire nc22034;
wire nc22035;
wire nc22036;
wire nc22037;
wire nc22038;
wire nc22039;
wire nc22040;
wire nc22041;
wire nc22042;
wire nc22043;
wire nc22044;
wire nc22045;
wire nc22046;
wire nc22047;
wire nc22048;
wire nc22049;
wire nc22050;
wire nc22051;
wire nc22052;
wire nc22053;
wire nc22054;
wire nc22055;
wire nc22056;
wire nc22057;
wire nc22058;
wire nc22059;
wire nc22060;
wire nc22061;
wire nc22062;
wire nc22063;
wire nc22064;
wire nc22065;
wire nc22066;
wire nc22067;
wire nc22068;
wire nc22069;
wire nc22070;
wire nc22071;
wire nc22072;
wire nc22073;
wire nc22074;
wire nc22075;
wire nc22076;
wire nc22077;
wire nc22078;
wire nc22079;
wire nc22080;
wire nc22081;
wire nc22082;
wire nc22083;
wire nc22084;
wire nc22085;
wire nc22086;
wire nc22087;
wire nc22088;
wire nc22089;
wire nc22090;
wire nc22091;
wire nc22092;
wire nc22093;
wire nc22094;
wire nc22095;
wire nc22096;
wire nc22097;
wire nc22098;
wire nc22099;
wire nc22100;
wire nc22101;
wire nc22102;
wire nc22103;
wire nc22104;
wire nc22105;
wire nc22106;
wire nc22107;
wire nc22108;
wire nc22109;
wire nc22110;
wire nc22111;
wire nc22112;
wire nc22113;
wire nc22114;
wire nc22115;
wire nc22116;
wire nc22117;
wire nc22118;
wire nc22119;
wire nc22120;
wire nc22121;
wire nc22122;
wire nc22123;
wire nc22124;
wire nc22125;
wire nc22126;
wire nc22127;
wire nc22128;
wire nc22129;
wire nc22130;
wire nc22131;
wire nc22132;
wire nc22133;
wire nc22134;
wire nc22135;
wire nc22136;
wire nc22137;
wire nc22138;
wire nc22139;
wire nc22140;
wire nc22141;
wire nc22142;
wire nc22143;
wire nc22144;
wire nc22145;
wire nc22146;
wire nc22147;
wire nc22148;
wire nc22149;
wire nc22150;
wire nc22151;
wire nc22152;
wire nc22153;
wire nc22154;
wire nc22155;
wire nc22156;
wire nc22157;
wire nc22158;
wire nc22159;
wire nc22160;
wire nc22161;
wire nc22162;
wire nc22163;
wire nc22164;
wire nc22165;
wire nc22166;
wire nc22167;
wire nc22168;
wire nc22169;
wire nc22170;
wire nc22171;
wire nc22172;
wire nc22173;
wire nc22174;
wire nc22175;
wire nc22176;
wire nc22177;
wire nc22178;
wire nc22179;
wire nc22180;
wire nc22181;
wire nc22182;
wire nc22183;
wire nc22184;
wire nc22185;
wire nc22186;
wire nc22187;
wire nc22188;
wire nc22189;
wire nc22190;
wire nc22191;
wire nc22192;
wire nc22193;
wire nc22194;
wire nc22195;
wire nc22196;
wire nc22197;
wire nc22198;
wire nc22199;
wire nc22200;
wire nc22201;
wire nc22202;
wire nc22203;
wire nc22204;
wire nc22205;
wire nc22206;
wire nc22207;
wire nc22208;
wire nc22209;
wire nc22210;
wire nc22211;
wire nc22212;
wire nc22213;
wire nc22214;
wire nc22215;
wire nc22216;
wire nc22217;
wire nc22218;
wire nc22219;
wire nc22220;
wire nc22221;
wire nc22222;
wire nc22223;
wire nc22224;
wire nc22225;
wire nc22226;
wire nc22227;
wire nc22228;
wire nc22229;
wire nc22230;
wire nc22231;
wire nc22232;
wire nc22233;
wire nc22234;
wire nc22235;
wire nc22236;
wire nc22237;
wire nc22238;
wire nc22239;
wire nc22240;
wire nc22241;
wire nc22242;
wire nc22243;
wire nc22244;
wire nc22245;
wire nc22246;
wire nc22247;
wire nc22248;
wire nc22249;
wire nc22250;
wire nc22251;
wire nc22252;
wire nc22253;
wire nc22254;
wire nc22255;
wire nc22256;
wire nc22257;
wire nc22258;
wire nc22259;
wire nc22260;
wire nc22261;
wire nc22262;
wire nc22263;
wire nc22264;
wire nc22265;
wire nc22266;
wire nc22267;
wire nc22268;
wire nc22269;
wire nc22270;
wire nc22271;
wire nc22272;
wire nc22273;
wire nc22274;
wire nc22275;
wire nc22276;
wire nc22277;
wire nc22278;
wire nc22279;
wire nc22280;
wire nc22281;
wire nc22282;
wire nc22283;
wire nc22284;
wire nc22285;
wire nc22286;
wire nc22287;
wire nc22288;
wire nc22289;
wire nc22290;
wire nc22291;
wire nc22292;
wire nc22293;
wire nc22294;
wire nc22295;
wire nc22296;
wire nc22297;
wire nc22298;
wire nc22299;
wire nc22300;
wire nc22301;
wire nc22302;
wire nc22303;
wire nc22304;
wire nc22305;
wire nc22306;
wire nc22307;
wire nc22308;
wire nc22309;
wire nc22310;
wire nc22311;
wire nc22312;
wire nc22313;
wire nc22314;
wire nc22315;
wire nc22316;
wire nc22317;
wire nc22318;
wire nc22319;
wire nc22320;
wire nc22321;
wire nc22322;
wire nc22323;
wire nc22324;
wire nc22325;
wire nc22326;
wire nc22327;
wire nc22328;
wire nc22329;
wire nc22330;
wire nc22331;
wire nc22332;
wire nc22333;
wire nc22334;
wire nc22335;
wire nc22336;
wire nc22337;
wire nc22338;
wire nc22339;
wire nc22340;
wire nc22341;
wire nc22342;
wire nc22343;
wire nc22344;
wire nc22345;
wire nc22346;
wire nc22347;
wire nc22348;
wire nc22349;
wire nc22350;
wire nc22351;
wire nc22352;
wire nc22353;
wire nc22354;
wire nc22355;
wire nc22356;
wire nc22357;
wire nc22358;
wire nc22359;
wire nc22360;
wire nc22361;
wire nc22362;
wire nc22363;
wire nc22364;
wire nc22365;
wire nc22366;
wire nc22367;
wire nc22368;
wire nc22369;
wire nc22370;
wire nc22371;
wire nc22372;
wire nc22373;
wire nc22374;
wire nc22375;
wire nc22376;
wire nc22377;
wire nc22378;
wire nc22379;
wire nc22380;
wire nc22381;
wire nc22382;
wire nc22383;
wire nc22384;
wire nc22385;
wire nc22386;
wire nc22387;
wire nc22388;
wire nc22389;
wire nc22390;
wire nc22391;
wire nc22392;
wire nc22393;
wire nc22394;
wire nc22395;
wire nc22396;
wire nc22397;
wire nc22398;
wire nc22399;
wire nc22400;
wire nc22401;
wire nc22402;
wire nc22403;
wire nc22404;
wire nc22405;
wire nc22406;
wire nc22407;
wire nc22408;
wire nc22409;
wire nc22410;
wire nc22411;
wire nc22412;
wire nc22413;
wire nc22414;
wire nc22415;
wire nc22416;
wire nc22417;
wire nc22418;
wire nc22419;
wire nc22420;
wire nc22421;
wire nc22422;
wire nc22423;
wire nc22424;
wire nc22425;
wire nc22426;
wire nc22427;
wire nc22428;
wire nc22429;
wire nc22430;
wire nc22431;
wire nc22432;
wire nc22433;
wire nc22434;
wire nc22435;
wire nc22436;
wire nc22437;
wire nc22438;
wire nc22439;
wire nc22440;
wire nc22441;
wire nc22442;
wire nc22443;
wire nc22444;
wire nc22445;
wire nc22446;
wire nc22447;
wire nc22448;
wire nc22449;
wire nc22450;
wire nc22451;
wire nc22452;
wire nc22453;
wire nc22454;
wire nc22455;
wire nc22456;
wire nc22457;
wire nc22458;
wire nc22459;
wire nc22460;
wire nc22461;
wire nc22462;
wire nc22463;
wire nc22464;
wire nc22465;
wire nc22466;
wire nc22467;
wire nc22468;
wire nc22469;
wire nc22470;
wire nc22471;
wire nc22472;
wire nc22473;
wire nc22474;
wire nc22475;
wire nc22476;
wire nc22477;
wire nc22478;
wire nc22479;
wire nc22480;
wire nc22481;
wire nc22482;
wire nc22483;
wire nc22484;
wire nc22485;
wire nc22486;
wire nc22487;
wire nc22488;
wire nc22489;
wire nc22490;
wire nc22491;
wire nc22492;
wire nc22493;
wire nc22494;
wire nc22495;
wire nc22496;
wire nc22497;
wire nc22498;
wire nc22499;
wire nc22500;
wire nc22501;
wire nc22502;
wire nc22503;
wire nc22504;
wire nc22505;
wire nc22506;
wire nc22507;
wire nc22508;
wire nc22509;
wire nc22510;
wire nc22511;
wire nc22512;
wire nc22513;
wire nc22514;
wire nc22515;
wire nc22516;
wire nc22517;
wire nc22518;
wire nc22519;
wire nc22520;
wire nc22521;
wire nc22522;
wire nc22523;
wire nc22524;
wire nc22525;
wire nc22526;
wire nc22527;
wire nc22528;
wire nc22529;
wire nc22530;
wire nc22531;
wire nc22532;
wire nc22533;
wire nc22534;
wire nc22535;
wire nc22536;
wire nc22537;
wire nc22538;
wire nc22539;
wire nc22540;
wire nc22541;
wire nc22542;
wire nc22543;
wire nc22544;
wire nc22545;
wire nc22546;
wire nc22547;
wire nc22548;
wire nc22549;
wire nc22550;
wire nc22551;
wire nc22552;
wire nc22553;
wire nc22554;
wire nc22555;
wire nc22556;
wire nc22557;
wire nc22558;
wire nc22559;
wire nc22560;
wire nc22561;
wire nc22562;
wire nc22563;
wire nc22564;
wire nc22565;
wire nc22566;
wire nc22567;
wire nc22568;
wire nc22569;
wire nc22570;
wire nc22571;
wire nc22572;
wire nc22573;
wire nc22574;
wire nc22575;
wire nc22576;
wire nc22577;
wire nc22578;
wire nc22579;
wire nc22580;
wire nc22581;
wire nc22582;
wire nc22583;
wire nc22584;
wire nc22585;
wire nc22586;
wire nc22587;
wire nc22588;
wire nc22589;
wire nc22590;
wire nc22591;
wire nc22592;
wire nc22593;
wire nc22594;
wire nc22595;
wire nc22596;
wire nc22597;
wire nc22598;
wire nc22599;
wire nc22600;
wire nc22601;
wire nc22602;
wire nc22603;
wire nc22604;
wire nc22605;
wire nc22606;
wire nc22607;
wire nc22608;
wire nc22609;
wire nc22610;
wire nc22611;
wire nc22612;
wire nc22613;
wire nc22614;
wire nc22615;
wire nc22616;
wire nc22617;
wire nc22618;
wire nc22619;
wire nc22620;
wire nc22621;
wire nc22622;
wire nc22623;
wire nc22624;
wire nc22625;
wire nc22626;
wire nc22627;
wire nc22628;
wire nc22629;
wire nc22630;
wire nc22631;
wire nc22632;
wire nc22633;
wire nc22634;
wire nc22635;
wire nc22636;
wire nc22637;
wire nc22638;
wire nc22639;
wire nc22640;
wire nc22641;
wire nc22642;
wire nc22643;
wire nc22644;
wire nc22645;
wire nc22646;
wire nc22647;
wire nc22648;
wire nc22649;
wire nc22650;
wire nc22651;
wire nc22652;
wire nc22653;
wire nc22654;
wire nc22655;
wire nc22656;
wire nc22657;
wire nc22658;
wire nc22659;
wire nc22660;
wire nc22661;
wire nc22662;
wire nc22663;
wire nc22664;
wire nc22665;
wire nc22666;
wire nc22667;
wire nc22668;
wire nc22669;
wire nc22670;
wire nc22671;
wire nc22672;
wire nc22673;
wire nc22674;
wire nc22675;
wire nc22676;
wire nc22677;
wire nc22678;
wire nc22679;
wire nc22680;
wire nc22681;
wire nc22682;
wire nc22683;
wire nc22684;
wire nc22685;
wire nc22686;
wire nc22687;
wire nc22688;
wire nc22689;
wire nc22690;
wire nc22691;
wire nc22692;
wire nc22693;
wire nc22694;
wire nc22695;
wire nc22696;
wire nc22697;
wire nc22698;
wire nc22699;
wire nc22700;
wire nc22701;
wire nc22702;
wire nc22703;
wire nc22704;
wire nc22705;
wire nc22706;
wire nc22707;
wire nc22708;
wire nc22709;
wire nc22710;
wire nc22711;
wire nc22712;
wire nc22713;
wire nc22714;
wire nc22715;
wire nc22716;
wire nc22717;
wire nc22718;
wire nc22719;
wire nc22720;
wire nc22721;
wire nc22722;
wire nc22723;
wire nc22724;
wire nc22725;
wire nc22726;
wire nc22727;
wire nc22728;
wire nc22729;
wire nc22730;
wire nc22731;
wire nc22732;
wire nc22733;
wire nc22734;
wire nc22735;
wire nc22736;
wire nc22737;
wire nc22738;
wire nc22739;
wire nc22740;
wire nc22741;
wire nc22742;
wire nc22743;
wire nc22744;
wire nc22745;
wire nc22746;
wire nc22747;
wire nc22748;
wire nc22749;
wire nc22750;
wire nc22751;
wire nc22752;
wire nc22753;
wire nc22754;
wire nc22755;
wire nc22756;
wire nc22757;
wire nc22758;
wire nc22759;
wire nc22760;
wire nc22761;
wire nc22762;
wire nc22763;
wire nc22764;
wire nc22765;
wire nc22766;
wire nc22767;
wire nc22768;
wire nc22769;
wire nc22770;
wire nc22771;
wire nc22772;
wire nc22773;
wire nc22774;
wire nc22775;
wire nc22776;
wire nc22777;
wire nc22778;
wire nc22779;
wire nc22780;
wire nc22781;
wire nc22782;
wire nc22783;
wire nc22784;
wire nc22785;
wire nc22786;
wire nc22787;
wire nc22788;
wire nc22789;
wire nc22790;
wire nc22791;
wire nc22792;
wire nc22793;
wire nc22794;
wire nc22795;
wire nc22796;
wire nc22797;
wire nc22798;
wire nc22799;
wire nc22800;
wire nc22801;
wire nc22802;
wire nc22803;
wire nc22804;
wire nc22805;
wire nc22806;
wire nc22807;
wire nc22808;
wire nc22809;
wire nc22810;
wire nc22811;
wire nc22812;
wire nc22813;
wire nc22814;
wire nc22815;
wire nc22816;
wire nc22817;
wire nc22818;
wire nc22819;
wire nc22820;
wire nc22821;
wire nc22822;
wire nc22823;
wire nc22824;
wire nc22825;
wire nc22826;
wire nc22827;
wire nc22828;
wire nc22829;
wire nc22830;
wire nc22831;
wire nc22832;
wire nc22833;
wire nc22834;
wire nc22835;
wire nc22836;
wire nc22837;
wire nc22838;
wire nc22839;
wire nc22840;
wire nc22841;
wire nc22842;
wire nc22843;
wire nc22844;
wire nc22845;
wire nc22846;
wire nc22847;
wire nc22848;
wire nc22849;
wire nc22850;
wire nc22851;
wire nc22852;
wire nc22853;
wire nc22854;
wire nc22855;
wire nc22856;
wire nc22857;
wire nc22858;
wire nc22859;
wire nc22860;
wire nc22861;
wire nc22862;
wire nc22863;
wire nc22864;
wire nc22865;
wire nc22866;
wire nc22867;
wire nc22868;
wire nc22869;
wire nc22870;
wire nc22871;
wire nc22872;
wire nc22873;
wire nc22874;
wire nc22875;
wire nc22876;
wire nc22877;
wire nc22878;
wire nc22879;
wire nc22880;
wire nc22881;
wire nc22882;
wire nc22883;
wire nc22884;
wire nc22885;
wire nc22886;
wire nc22887;
wire nc22888;
wire nc22889;
wire nc22890;
wire nc22891;
wire nc22892;
wire nc22893;
wire nc22894;
wire nc22895;
wire nc22896;
wire nc22897;
wire nc22898;
wire nc22899;
wire nc22900;
wire nc22901;
wire nc22902;
wire nc22903;
wire nc22904;
wire nc22905;
wire nc22906;
wire nc22907;
wire nc22908;
wire nc22909;
wire nc22910;
wire nc22911;
wire nc22912;
wire nc22913;
wire nc22914;
wire nc22915;
wire nc22916;
wire nc22917;
wire nc22918;
wire nc22919;
wire nc22920;
wire nc22921;
wire nc22922;
wire nc22923;
wire nc22924;
wire nc22925;
wire nc22926;
wire nc22927;
wire nc22928;
wire nc22929;
wire nc22930;
wire nc22931;
wire nc22932;
wire nc22933;
wire nc22934;
wire nc22935;
wire nc22936;
wire nc22937;
wire nc22938;
wire nc22939;
wire nc22940;
wire nc22941;
wire nc22942;
wire nc22943;
wire nc22944;
wire nc22945;
wire nc22946;
wire nc22947;
wire nc22948;
wire nc22949;
wire nc22950;
wire nc22951;
wire nc22952;
wire nc22953;
wire nc22954;
wire nc22955;
wire nc22956;
wire nc22957;
wire nc22958;
wire nc22959;
wire nc22960;
wire nc22961;
wire nc22962;
wire nc22963;
wire nc22964;
wire nc22965;
wire nc22966;
wire nc22967;
wire nc22968;
wire nc22969;
wire nc22970;
wire nc22971;
wire nc22972;
wire nc22973;
wire nc22974;
wire nc22975;
wire nc22976;
wire nc22977;
wire nc22978;
wire nc22979;
wire nc22980;
wire nc22981;
wire nc22982;
wire nc22983;
wire nc22984;
wire nc22985;
wire nc22986;
wire nc22987;
wire nc22988;
wire nc22989;
wire nc22990;
wire nc22991;
wire nc22992;
wire nc22993;
wire nc22994;
wire nc22995;
wire nc22996;
wire nc22997;
wire nc22998;
wire nc22999;
wire nc23000;
wire nc23001;
wire nc23002;
wire nc23003;
wire nc23004;
wire nc23005;
wire nc23006;
wire nc23007;
wire nc23008;
wire nc23009;
wire nc23010;
wire nc23011;
wire nc23012;
wire nc23013;
wire nc23014;
wire nc23015;
wire nc23016;
wire nc23017;
wire nc23018;
wire nc23019;
wire nc23020;
wire nc23021;
wire nc23022;
wire nc23023;
wire nc23024;
wire nc23025;
wire nc23026;
wire nc23027;
wire nc23028;
wire nc23029;
wire nc23030;
wire nc23031;
wire nc23032;
wire nc23033;
wire nc23034;
wire nc23035;
wire nc23036;
wire nc23037;
wire nc23038;
wire nc23039;
wire nc23040;
wire nc23041;
wire nc23042;
wire nc23043;
wire nc23044;
wire nc23045;
wire nc23046;
wire nc23047;
wire nc23048;
wire nc23049;
wire nc23050;
wire nc23051;
wire nc23052;
wire nc23053;
wire nc23054;
wire nc23055;
wire nc23056;
wire nc23057;
wire nc23058;
wire nc23059;
wire nc23060;
wire nc23061;
wire nc23062;
wire nc23063;
wire nc23064;
wire nc23065;
wire nc23066;
wire nc23067;
wire nc23068;
wire nc23069;
wire nc23070;
wire nc23071;
wire nc23072;
wire nc23073;
wire nc23074;
wire nc23075;
wire nc23076;
wire nc23077;
wire nc23078;
wire nc23079;
wire nc23080;
wire nc23081;
wire nc23082;
wire nc23083;
wire nc23084;
wire nc23085;
wire nc23086;
wire nc23087;
wire nc23088;
wire nc23089;
wire nc23090;
wire nc23091;
wire nc23092;
wire nc23093;
wire nc23094;
wire nc23095;
wire nc23096;
wire nc23097;
wire nc23098;
wire nc23099;
wire nc23100;
wire nc23101;
wire nc23102;
wire nc23103;
wire nc23104;
wire nc23105;
wire nc23106;
wire nc23107;
wire nc23108;
wire nc23109;
wire nc23110;
wire nc23111;
wire nc23112;
wire nc23113;
wire nc23114;
wire nc23115;
wire nc23116;
wire nc23117;
wire nc23118;
wire nc23119;
wire nc23120;
wire nc23121;
wire nc23122;
wire nc23123;
wire nc23124;
wire nc23125;
wire nc23126;
wire nc23127;
wire nc23128;
wire nc23129;
wire nc23130;
wire nc23131;
wire nc23132;
wire nc23133;
wire nc23134;
wire nc23135;
wire nc23136;
wire nc23137;
wire nc23138;
wire nc23139;
wire nc23140;
wire nc23141;
wire nc23142;
wire nc23143;
wire nc23144;
wire nc23145;
wire nc23146;
wire nc23147;
wire nc23148;
wire nc23149;
wire nc23150;
wire nc23151;
wire nc23152;
wire nc23153;
wire nc23154;
wire nc23155;
wire nc23156;
wire nc23157;
wire nc23158;
wire nc23159;
wire nc23160;
wire nc23161;
wire nc23162;
wire nc23163;
wire nc23164;
wire nc23165;
wire nc23166;
wire nc23167;
wire nc23168;
wire nc23169;
wire nc23170;
wire nc23171;
wire nc23172;
wire nc23173;
wire nc23174;
wire nc23175;
wire nc23176;
wire nc23177;
wire nc23178;
wire nc23179;
wire nc23180;
wire nc23181;
wire nc23182;
wire nc23183;
wire nc23184;
wire nc23185;
wire nc23186;
wire nc23187;
wire nc23188;
wire nc23189;
wire nc23190;
wire nc23191;
wire nc23192;
wire nc23193;
wire nc23194;
wire nc23195;
wire nc23196;
wire nc23197;
wire nc23198;
wire nc23199;
wire nc23200;
wire nc23201;
wire nc23202;
wire nc23203;
wire nc23204;
wire nc23205;
wire nc23206;
wire nc23207;
wire nc23208;
wire nc23209;
wire nc23210;
wire nc23211;
wire nc23212;
wire nc23213;
wire nc23214;
wire nc23215;
wire nc23216;
wire nc23217;
wire nc23218;
wire nc23219;
wire nc23220;
wire nc23221;
wire nc23222;
wire nc23223;
wire nc23224;
wire nc23225;
wire nc23226;
wire nc23227;
wire nc23228;
wire nc23229;
wire nc23230;
wire nc23231;
wire nc23232;
wire nc23233;
wire nc23234;
wire nc23235;
wire nc23236;
wire nc23237;
wire nc23238;
wire nc23239;
wire nc23240;
wire nc23241;
wire nc23242;
wire nc23243;
wire nc23244;
wire nc23245;
wire nc23246;
wire nc23247;
wire nc23248;
wire nc23249;
wire nc23250;
wire nc23251;
wire nc23252;
wire nc23253;
wire nc23254;
wire nc23255;
wire nc23256;
wire nc23257;
wire nc23258;
wire nc23259;
wire nc23260;
wire nc23261;
wire nc23262;
wire nc23263;
wire nc23264;
wire nc23265;
wire nc23266;
wire nc23267;
wire nc23268;
wire nc23269;
wire nc23270;
wire nc23271;
wire nc23272;
wire nc23273;
wire nc23274;
wire nc23275;
wire nc23276;
wire nc23277;
wire nc23278;
wire nc23279;
wire nc23280;
wire nc23281;
wire nc23282;
wire nc23283;
wire nc23284;
wire nc23285;
wire nc23286;
wire nc23287;
wire nc23288;
wire nc23289;
wire nc23290;
wire nc23291;
wire nc23292;
wire nc23293;
wire nc23294;
wire nc23295;
wire nc23296;
wire nc23297;
wire nc23298;
wire nc23299;
wire nc23300;
wire nc23301;
wire nc23302;
wire nc23303;
wire nc23304;
wire nc23305;
wire nc23306;
wire nc23307;
wire nc23308;
wire nc23309;
wire nc23310;
wire nc23311;
wire nc23312;
wire nc23313;
wire nc23314;
wire nc23315;
wire nc23316;
wire nc23317;
wire nc23318;
wire nc23319;
wire nc23320;
wire nc23321;
wire nc23322;
wire nc23323;
wire nc23324;
wire nc23325;
wire nc23326;
wire nc23327;
wire nc23328;
wire nc23329;
wire nc23330;
wire nc23331;
wire nc23332;
wire nc23333;
wire nc23334;
wire nc23335;
wire nc23336;
wire nc23337;
wire nc23338;
wire nc23339;
wire nc23340;
wire nc23341;
wire nc23342;
wire nc23343;
wire nc23344;
wire nc23345;
wire nc23346;
wire nc23347;
wire nc23348;
wire nc23349;
wire nc23350;
wire nc23351;
wire nc23352;
wire nc23353;
wire nc23354;
wire nc23355;
wire nc23356;
wire nc23357;
wire nc23358;
wire nc23359;
wire nc23360;
wire nc23361;
wire nc23362;
wire nc23363;
wire nc23364;
wire nc23365;
wire nc23366;
wire nc23367;
wire nc23368;
wire nc23369;
wire nc23370;
wire nc23371;
wire nc23372;
wire nc23373;
wire nc23374;
wire nc23375;
wire nc23376;
wire nc23377;
wire nc23378;
wire nc23379;
wire nc23380;
wire nc23381;
wire nc23382;
wire nc23383;
wire nc23384;
wire nc23385;
wire nc23386;
wire nc23387;
wire nc23388;
wire nc23389;
wire nc23390;
wire nc23391;
wire nc23392;
wire nc23393;
wire nc23394;
wire nc23395;
wire nc23396;
wire nc23397;
wire nc23398;
wire nc23399;
wire nc23400;
wire nc23401;
wire nc23402;
wire nc23403;
wire nc23404;
wire nc23405;
wire nc23406;
wire nc23407;
wire nc23408;
wire nc23409;
wire nc23410;
wire nc23411;
wire nc23412;
wire nc23413;
wire nc23414;
wire nc23415;
wire nc23416;
wire nc23417;
wire nc23418;
wire nc23419;
wire nc23420;
wire nc23421;
wire nc23422;
wire nc23423;
wire nc23424;
wire nc23425;
wire nc23426;
wire nc23427;
wire nc23428;
wire nc23429;
wire nc23430;
wire nc23431;
wire nc23432;
wire nc23433;
wire nc23434;
wire nc23435;
wire nc23436;
wire nc23437;
wire nc23438;
wire nc23439;
wire nc23440;
wire nc23441;
wire nc23442;
wire nc23443;
wire nc23444;
wire nc23445;
wire nc23446;
wire nc23447;
wire nc23448;
wire nc23449;
wire nc23450;
wire nc23451;
wire nc23452;
wire nc23453;
wire nc23454;
wire nc23455;
wire nc23456;
wire nc23457;
wire nc23458;
wire nc23459;
wire nc23460;
wire nc23461;
wire nc23462;
wire nc23463;
wire nc23464;
wire nc23465;
wire nc23466;
wire nc23467;
wire nc23468;
wire nc23469;
wire nc23470;
wire nc23471;
wire nc23472;
wire nc23473;
wire nc23474;
wire nc23475;
wire nc23476;
wire nc23477;
wire nc23478;
wire nc23479;
wire nc23480;
wire nc23481;
wire nc23482;
wire nc23483;
wire nc23484;
wire nc23485;
wire nc23486;
wire nc23487;
wire nc23488;
wire nc23489;
wire nc23490;
wire nc23491;
wire nc23492;
wire nc23493;
wire nc23494;
wire nc23495;
wire nc23496;
wire nc23497;
wire nc23498;
wire nc23499;
wire nc23500;
wire nc23501;
wire nc23502;
wire nc23503;
wire nc23504;
wire nc23505;
wire nc23506;
wire nc23507;
wire nc23508;
wire nc23509;
wire nc23510;
wire nc23511;
wire nc23512;
wire nc23513;
wire nc23514;
wire nc23515;
wire nc23516;
wire nc23517;
wire nc23518;
wire nc23519;
wire nc23520;
wire nc23521;
wire nc23522;
wire nc23523;
wire nc23524;
wire nc23525;
wire nc23526;
wire nc23527;
wire nc23528;
wire nc23529;
wire nc23530;
wire nc23531;
wire nc23532;
wire nc23533;
wire nc23534;
wire nc23535;
wire nc23536;
wire nc23537;
wire nc23538;
wire nc23539;
wire nc23540;
wire nc23541;
wire nc23542;
wire nc23543;
wire nc23544;
wire nc23545;
wire nc23546;
wire nc23547;
wire nc23548;
wire nc23549;
wire nc23550;
wire nc23551;
wire nc23552;
wire nc23553;
wire nc23554;
wire nc23555;
wire nc23556;
wire nc23557;
wire nc23558;
wire nc23559;
wire nc23560;
wire nc23561;
wire nc23562;
wire nc23563;
wire nc23564;
wire nc23565;
wire nc23566;
wire nc23567;
wire nc23568;
wire nc23569;
wire nc23570;
wire nc23571;
wire nc23572;
wire nc23573;
wire nc23574;
wire nc23575;
wire nc23576;
wire nc23577;
wire nc23578;
wire nc23579;
wire nc23580;
wire nc23581;
wire nc23582;
wire nc23583;
wire nc23584;
wire nc23585;
wire nc23586;
wire nc23587;
wire nc23588;
wire nc23589;
wire nc23590;
wire nc23591;
wire nc23592;
wire nc23593;
wire nc23594;
wire nc23595;
wire nc23596;
wire nc23597;
wire nc23598;
wire nc23599;
wire nc23600;
wire nc23601;
wire nc23602;
wire nc23603;
wire nc23604;
wire nc23605;
wire nc23606;
wire nc23607;
wire nc23608;
wire nc23609;
wire nc23610;
wire nc23611;
wire nc23612;
wire nc23613;
wire nc23614;
wire nc23615;
wire nc23616;
wire nc23617;
wire nc23618;
wire nc23619;
wire nc23620;
wire nc23621;
wire nc23622;
wire nc23623;
wire nc23624;
wire nc23625;
wire nc23626;
wire nc23627;
wire nc23628;
wire nc23629;
wire nc23630;
wire nc23631;
wire nc23632;
wire nc23633;
wire nc23634;
wire nc23635;
wire nc23636;
wire nc23637;
wire nc23638;
wire nc23639;
wire nc23640;
wire nc23641;
wire nc23642;
wire nc23643;
wire nc23644;
wire nc23645;
wire nc23646;
wire nc23647;
wire nc23648;
wire nc23649;
wire nc23650;
wire nc23651;
wire nc23652;
wire nc23653;
wire nc23654;
wire nc23655;
wire nc23656;
wire nc23657;
wire nc23658;
wire nc23659;
wire nc23660;
wire nc23661;
wire nc23662;
wire nc23663;
wire nc23664;
wire nc23665;
wire nc23666;
wire nc23667;
wire nc23668;
wire nc23669;
wire nc23670;
wire nc23671;
wire nc23672;
wire nc23673;
wire nc23674;
wire nc23675;
wire nc23676;
wire nc23677;
wire nc23678;
wire nc23679;
wire nc23680;
wire nc23681;
wire nc23682;
wire nc23683;
wire nc23684;
wire nc23685;
wire nc23686;
wire nc23687;
wire nc23688;
wire nc23689;
wire nc23690;
wire nc23691;
wire nc23692;
wire nc23693;
wire nc23694;
wire nc23695;
wire nc23696;
wire nc23697;
wire nc23698;
wire nc23699;
wire nc23700;
wire nc23701;
wire nc23702;
wire nc23703;
wire nc23704;
wire nc23705;
wire nc23706;
wire nc23707;
wire nc23708;
wire nc23709;
wire nc23710;
wire nc23711;
wire nc23712;
wire nc23713;
wire nc23714;
wire nc23715;
wire nc23716;
wire nc23717;
wire nc23718;
wire nc23719;
wire nc23720;
wire nc23721;
wire nc23722;
wire nc23723;
wire nc23724;
wire nc23725;
wire nc23726;
wire nc23727;
wire nc23728;
wire nc23729;
wire nc23730;
wire nc23731;
wire nc23732;
wire nc23733;
wire nc23734;
wire nc23735;
wire nc23736;
wire nc23737;
wire nc23738;
wire nc23739;
wire nc23740;
wire nc23741;
wire nc23742;
wire nc23743;
wire nc23744;
wire nc23745;
wire nc23746;
wire nc23747;
wire nc23748;
wire nc23749;
wire nc23750;
wire nc23751;
wire nc23752;
wire nc23753;
wire nc23754;
wire nc23755;
wire nc23756;
wire nc23757;
wire nc23758;
wire nc23759;
wire nc23760;
wire nc23761;
wire nc23762;
wire nc23763;
wire nc23764;
wire nc23765;
wire nc23766;
wire nc23767;
wire nc23768;
wire nc23769;
wire nc23770;
wire nc23771;
wire nc23772;
wire nc23773;
wire nc23774;
wire nc23775;
wire nc23776;
wire nc23777;
wire nc23778;
wire nc23779;
wire nc23780;
wire nc23781;
wire nc23782;
wire nc23783;
wire nc23784;
wire nc23785;
wire nc23786;
wire nc23787;
wire nc23788;
wire nc23789;
wire nc23790;
wire nc23791;
wire nc23792;
wire nc23793;
wire nc23794;
wire nc23795;
wire nc23796;
wire nc23797;
wire nc23798;
wire nc23799;
wire nc23800;
wire nc23801;
wire nc23802;
wire nc23803;
wire nc23804;
wire nc23805;
wire nc23806;
wire nc23807;
wire nc23808;
wire nc23809;
wire nc23810;
wire nc23811;
wire nc23812;
wire nc23813;
wire nc23814;
wire nc23815;
wire nc23816;
wire nc23817;
wire nc23818;
wire nc23819;
wire nc23820;
wire nc23821;
wire nc23822;
wire nc23823;
wire nc23824;
wire nc23825;
wire nc23826;
wire nc23827;
wire nc23828;
wire nc23829;
wire nc23830;
wire nc23831;
wire nc23832;
wire nc23833;
wire nc23834;
wire nc23835;
wire nc23836;
wire nc23837;
wire nc23838;
wire nc23839;
wire nc23840;
wire nc23841;
wire nc23842;
wire nc23843;
wire nc23844;
wire nc23845;
wire nc23846;
wire nc23847;
wire nc23848;
wire nc23849;
wire nc23850;
wire nc23851;
wire nc23852;
wire nc23853;
wire nc23854;
wire nc23855;
wire nc23856;
wire nc23857;
wire nc23858;
wire nc23859;
wire nc23860;
wire nc23861;
wire nc23862;
wire nc23863;
wire nc23864;
wire nc23865;
wire nc23866;
wire nc23867;
wire nc23868;
wire nc23869;
wire nc23870;
wire nc23871;
wire nc23872;
wire nc23873;
wire nc23874;
wire nc23875;
wire nc23876;
wire nc23877;
wire nc23878;
wire nc23879;
wire nc23880;
wire nc23881;
wire nc23882;
wire nc23883;
wire nc23884;
wire nc23885;
wire nc23886;
wire nc23887;
wire nc23888;
wire nc23889;
wire nc23890;
wire nc23891;
wire nc23892;
wire nc23893;
wire nc23894;
wire nc23895;
wire nc23896;
wire nc23897;
wire nc23898;
wire nc23899;
wire nc23900;
wire nc23901;
wire nc23902;
wire nc23903;
wire nc23904;
wire nc23905;
wire nc23906;
wire nc23907;
wire nc23908;
wire nc23909;
wire nc23910;
wire nc23911;
wire nc23912;
wire nc23913;
wire nc23914;
wire nc23915;
wire nc23916;
wire nc23917;
wire nc23918;
wire nc23919;
wire nc23920;
wire nc23921;
wire nc23922;
wire nc23923;
wire nc23924;
wire nc23925;
wire nc23926;
wire nc23927;
wire nc23928;
wire nc23929;
wire nc23930;
wire nc23931;
wire nc23932;
wire nc23933;
wire nc23934;
wire nc23935;
wire nc23936;
wire nc23937;
wire nc23938;
wire nc23939;
wire nc23940;
wire nc23941;
wire nc23942;
wire nc23943;
wire nc23944;
wire nc23945;
wire nc23946;
wire nc23947;
wire nc23948;
wire nc23949;
wire nc23950;
wire nc23951;
wire nc23952;
wire nc23953;
wire nc23954;
wire nc23955;
wire nc23956;
wire nc23957;
wire nc23958;
wire nc23959;
wire nc23960;
wire nc23961;
wire nc23962;
wire nc23963;
wire nc23964;
wire nc23965;
wire nc23966;
wire nc23967;
wire nc23968;
wire nc23969;
wire nc23970;
wire nc23971;
wire nc23972;
wire nc23973;
wire nc23974;
wire nc23975;
wire nc23976;
wire nc23977;
wire nc23978;
wire nc23979;
wire nc23980;
wire nc23981;
wire nc23982;
wire nc23983;
wire nc23984;
wire nc23985;
wire nc23986;
wire nc23987;
wire nc23988;
wire nc23989;
wire nc23990;
wire nc23991;
wire nc23992;
wire nc23993;
wire nc23994;
wire nc23995;
wire nc23996;
wire nc23997;
wire nc23998;
wire nc23999;
wire nc24000;
wire nc24001;
wire nc24002;
wire nc24003;
wire nc24004;
wire nc24005;
wire nc24006;
wire nc24007;
wire nc24008;
wire nc24009;
wire nc24010;
wire nc24011;
wire nc24012;
wire nc24013;
wire nc24014;
wire nc24015;
wire nc24016;
wire nc24017;
wire nc24018;
wire nc24019;
wire nc24020;
wire nc24021;
wire nc24022;
wire nc24023;
wire nc24024;
wire nc24025;
wire nc24026;
wire nc24027;
wire nc24028;
wire nc24029;
wire nc24030;
wire nc24031;
wire nc24032;
wire nc24033;
wire nc24034;
wire nc24035;
wire nc24036;
wire nc24037;
wire nc24038;
wire nc24039;
wire nc24040;
wire nc24041;
wire nc24042;
wire nc24043;
wire nc24044;
wire nc24045;
wire nc24046;
wire nc24047;
wire nc24048;
wire nc24049;
wire nc24050;
wire nc24051;
wire nc24052;
wire nc24053;
wire nc24054;
wire nc24055;
wire nc24056;
wire nc24057;
wire nc24058;
wire nc24059;
wire nc24060;
wire nc24061;
wire nc24062;
wire nc24063;
wire nc24064;
wire nc24065;
wire nc24066;
wire nc24067;
wire nc24068;
wire nc24069;
wire nc24070;
wire nc24071;
wire nc24072;
wire nc24073;
wire nc24074;
wire nc24075;
wire nc24076;
wire nc24077;
wire nc24078;
wire nc24079;
wire nc24080;
wire nc24081;
wire nc24082;
wire nc24083;
wire nc24084;
wire nc24085;
wire nc24086;
wire nc24087;
wire nc24088;
wire nc24089;
wire nc24090;
wire nc24091;
wire nc24092;
wire nc24093;
wire nc24094;
wire nc24095;
wire nc24096;
wire nc24097;
wire nc24098;
wire nc24099;
wire nc24100;
wire nc24101;
wire nc24102;
wire nc24103;
wire nc24104;
wire nc24105;
wire nc24106;
wire nc24107;
wire nc24108;
wire nc24109;
wire nc24110;
wire nc24111;
wire nc24112;
wire nc24113;
wire nc24114;
wire nc24115;
wire nc24116;
wire nc24117;
wire nc24118;
wire nc24119;
wire nc24120;
wire nc24121;
wire nc24122;
wire nc24123;
wire nc24124;
wire nc24125;
wire nc24126;
wire nc24127;
wire nc24128;
wire nc24129;
wire nc24130;
wire nc24131;
wire nc24132;
wire nc24133;
wire nc24134;
wire nc24135;
wire nc24136;
wire nc24137;
wire nc24138;
wire nc24139;
wire nc24140;
wire nc24141;
wire nc24142;
wire nc24143;
wire nc24144;
wire nc24145;
wire nc24146;
wire nc24147;
wire nc24148;
wire nc24149;
wire nc24150;
wire nc24151;
wire nc24152;
wire nc24153;
wire nc24154;
wire nc24155;
wire nc24156;
wire nc24157;
wire nc24158;
wire nc24159;
wire nc24160;
wire nc24161;
wire nc24162;
wire nc24163;
wire nc24164;
wire nc24165;
wire nc24166;
wire nc24167;
wire nc24168;
wire nc24169;
wire nc24170;
wire nc24171;
wire nc24172;
wire nc24173;
wire nc24174;
wire nc24175;
wire nc24176;
wire nc24177;
wire nc24178;
wire nc24179;
wire nc24180;
wire nc24181;
wire nc24182;
wire nc24183;
wire nc24184;
wire nc24185;
wire nc24186;
wire nc24187;
wire nc24188;
wire nc24189;
wire nc24190;
wire nc24191;
wire nc24192;
wire nc24193;
wire nc24194;
wire nc24195;
wire nc24196;
wire nc24197;
wire nc24198;
wire nc24199;
wire nc24200;
wire nc24201;
wire nc24202;
wire nc24203;
wire nc24204;
wire nc24205;
wire nc24206;
wire nc24207;
wire nc24208;
wire nc24209;
wire nc24210;
wire nc24211;
wire nc24212;
wire nc24213;
wire nc24214;
wire nc24215;
wire nc24216;
wire nc24217;
wire nc24218;
wire nc24219;
wire nc24220;
wire nc24221;
wire nc24222;
wire nc24223;
wire nc24224;
wire nc24225;
wire nc24226;
wire nc24227;
wire nc24228;
wire nc24229;
wire nc24230;
wire nc24231;
wire nc24232;
wire nc24233;
wire nc24234;
wire nc24235;
wire nc24236;
wire nc24237;
wire nc24238;
wire nc24239;
wire nc24240;
wire nc24241;
wire nc24242;
wire nc24243;
wire nc24244;
wire nc24245;
wire nc24246;
wire nc24247;
wire nc24248;
wire nc24249;
wire nc24250;
wire nc24251;
wire nc24252;
wire nc24253;
wire nc24254;
wire nc24255;
wire nc24256;
wire nc24257;
wire nc24258;
wire nc24259;
wire nc24260;
wire nc24261;
wire nc24262;
wire nc24263;
wire nc24264;
wire nc24265;
wire nc24266;
wire nc24267;
wire nc24268;
wire nc24269;
wire nc24270;
wire nc24271;
wire nc24272;
wire nc24273;
wire nc24274;
wire nc24275;
wire nc24276;
wire nc24277;
wire nc24278;
wire nc24279;
wire nc24280;
wire nc24281;
wire nc24282;
wire nc24283;
wire nc24284;
wire nc24285;
wire nc24286;
wire nc24287;
wire nc24288;
wire nc24289;
wire nc24290;
wire nc24291;
wire nc24292;
wire nc24293;
wire nc24294;
wire nc24295;
wire nc24296;
wire nc24297;
wire nc24298;
wire nc24299;
wire nc24300;
wire nc24301;
wire nc24302;
wire nc24303;
wire nc24304;
wire nc24305;
wire nc24306;
wire nc24307;
wire nc24308;
wire nc24309;
wire nc24310;
wire nc24311;
wire nc24312;
wire nc24313;
wire nc24314;
wire nc24315;
wire nc24316;
wire nc24317;
wire nc24318;
wire nc24319;
wire nc24320;
wire nc24321;
wire nc24322;
wire nc24323;
wire nc24324;
wire nc24325;
wire nc24326;
wire nc24327;
wire nc24328;
wire nc24329;
wire nc24330;
wire nc24331;
wire nc24332;
wire nc24333;
wire nc24334;
wire nc24335;
wire nc24336;
wire nc24337;
wire nc24338;
wire nc24339;
wire nc24340;
wire nc24341;
wire nc24342;
wire nc24343;
wire nc24344;
wire nc24345;
wire nc24346;
wire nc24347;
wire nc24348;
wire nc24349;
wire nc24350;
wire nc24351;
wire nc24352;
wire nc24353;
wire nc24354;
wire nc24355;
wire nc24356;
wire nc24357;
wire nc24358;
wire nc24359;
wire nc24360;
wire nc24361;
wire nc24362;
wire nc24363;
wire nc24364;
wire nc24365;
wire nc24366;
wire nc24367;
wire nc24368;
wire nc24369;
wire nc24370;
wire nc24371;
wire nc24372;
wire nc24373;
wire nc24374;
wire nc24375;
wire nc24376;
wire nc24377;
wire nc24378;
wire nc24379;
wire nc24380;
wire nc24381;
wire nc24382;
wire nc24383;
wire nc24384;
wire nc24385;
wire nc24386;
wire nc24387;
wire nc24388;
wire nc24389;
wire nc24390;
wire nc24391;
wire nc24392;
wire nc24393;
wire nc24394;
wire nc24395;
wire nc24396;
wire nc24397;
wire nc24398;
wire nc24399;
wire nc24400;
wire nc24401;
wire nc24402;
wire nc24403;
wire nc24404;
wire nc24405;
wire nc24406;
wire nc24407;
wire nc24408;
wire nc24409;
wire nc24410;
wire nc24411;
wire nc24412;
wire nc24413;
wire nc24414;
wire nc24415;
wire nc24416;
wire nc24417;
wire nc24418;
wire nc24419;
wire nc24420;
wire nc24421;
wire nc24422;
wire nc24423;
wire nc24424;
wire nc24425;
wire nc24426;
wire nc24427;
wire nc24428;
wire nc24429;
wire nc24430;
wire nc24431;
wire nc24432;
wire nc24433;
wire nc24434;
wire nc24435;
wire nc24436;
wire nc24437;
wire nc24438;
wire nc24439;
wire nc24440;
wire nc24441;
wire nc24442;
wire nc24443;
wire nc24444;
wire nc24445;
wire nc24446;
wire nc24447;
wire nc24448;
wire nc24449;
wire nc24450;
wire nc24451;
wire nc24452;
wire nc24453;
wire nc24454;
wire nc24455;
wire nc24456;
wire nc24457;
wire nc24458;
wire nc24459;
wire nc24460;
wire nc24461;
wire nc24462;
wire nc24463;
wire nc24464;
wire nc24465;
wire nc24466;
wire nc24467;
wire nc24468;
wire nc24469;
wire nc24470;
wire nc24471;
wire nc24472;
wire nc24473;
wire nc24474;
wire nc24475;
wire nc24476;
wire nc24477;
wire nc24478;
wire nc24479;
wire nc24480;
wire nc24481;
wire nc24482;
wire nc24483;
wire nc24484;
wire nc24485;
wire nc24486;
wire nc24487;
wire nc24488;
wire nc24489;
wire nc24490;
wire nc24491;
wire nc24492;
wire nc24493;
wire nc24494;
wire nc24495;
wire nc24496;
wire nc24497;
wire nc24498;
wire nc24499;
wire nc24500;
wire nc24501;
wire nc24502;
wire nc24503;
wire nc24504;
wire nc24505;
wire nc24506;
wire nc24507;
wire nc24508;
wire nc24509;
wire nc24510;
wire nc24511;
wire nc24512;
wire nc24513;
wire nc24514;
wire nc24515;
wire nc24516;
wire nc24517;
wire nc24518;
wire nc24519;
wire nc24520;
wire nc24521;
wire nc24522;
wire nc24523;
wire nc24524;
wire nc24525;
wire nc24526;
wire nc24527;
wire nc24528;
wire nc24529;
wire nc24530;
wire nc24531;
wire nc24532;
wire nc24533;
wire nc24534;
wire nc24535;
wire nc24536;
wire nc24537;
wire nc24538;
wire nc24539;
wire nc24540;
wire nc24541;
wire nc24542;
wire nc24543;
wire nc24544;
wire nc24545;
wire nc24546;
wire nc24547;
wire nc24548;
wire nc24549;
wire nc24550;
wire nc24551;
wire nc24552;
wire nc24553;
wire nc24554;
wire nc24555;
wire nc24556;
wire nc24557;
wire nc24558;
wire nc24559;
wire nc24560;
wire nc24561;
wire nc24562;
wire nc24563;
wire nc24564;
wire nc24565;
wire nc24566;
wire nc24567;
wire nc24568;
wire nc24569;
wire nc24570;
wire nc24571;
wire nc24572;
wire nc24573;
wire nc24574;
wire nc24575;
wire nc24576;
wire nc24577;
wire nc24578;
wire nc24579;
wire nc24580;
wire nc24581;
wire nc24582;
wire nc24583;
wire nc24584;
wire nc24585;
wire nc24586;
wire nc24587;
wire nc24588;
wire nc24589;
wire nc24590;
wire nc24591;
wire nc24592;
wire nc24593;
wire nc24594;
wire nc24595;
wire nc24596;
wire nc24597;
wire nc24598;
wire nc24599;
wire nc24600;
wire nc24601;
wire nc24602;
wire nc24603;
wire nc24604;
wire nc24605;
wire nc24606;
wire nc24607;
wire nc24608;
wire nc24609;
wire nc24610;
wire nc24611;
wire nc24612;
wire nc24613;
wire nc24614;
wire nc24615;
wire nc24616;
wire nc24617;
wire nc24618;
wire nc24619;
wire nc24620;
wire nc24621;
wire nc24622;
wire nc24623;
wire nc24624;
wire nc24625;
wire nc24626;
wire nc24627;
wire nc24628;
wire nc24629;
wire nc24630;
wire nc24631;
wire nc24632;
wire nc24633;
wire nc24634;
wire nc24635;
wire nc24636;
wire nc24637;
wire nc24638;
wire nc24639;
wire nc24640;
wire nc24641;
wire nc24642;
wire nc24643;
wire nc24644;
wire nc24645;
wire nc24646;
wire nc24647;
wire nc24648;
wire nc24649;
wire nc24650;
wire nc24651;
wire nc24652;
wire nc24653;
wire nc24654;
wire nc24655;
wire nc24656;
wire nc24657;
wire nc24658;
wire nc24659;
wire nc24660;
wire nc24661;
wire nc24662;
wire nc24663;
wire nc24664;
wire nc24665;
wire nc24666;
wire nc24667;
wire nc24668;
wire nc24669;
wire nc24670;
wire nc24671;
wire nc24672;
wire nc24673;
wire nc24674;
wire nc24675;
wire nc24676;
wire nc24677;
wire nc24678;
wire nc24679;
wire nc24680;
wire nc24681;
wire nc24682;
wire nc24683;
wire nc24684;
wire nc24685;
wire nc24686;
wire nc24687;
wire nc24688;
wire nc24689;
wire nc24690;
wire nc24691;
wire nc24692;
wire nc24693;
wire nc24694;
wire nc24695;
wire nc24696;
wire nc24697;
wire nc24698;
wire nc24699;
wire nc24700;
wire nc24701;
wire nc24702;
wire nc24703;
wire nc24704;
wire nc24705;
wire nc24706;
wire nc24707;
wire nc24708;
wire nc24709;
wire nc24710;
wire nc24711;
wire nc24712;
wire nc24713;
wire nc24714;
wire nc24715;
wire nc24716;
wire nc24717;
wire nc24718;
wire nc24719;
wire nc24720;
wire nc24721;
wire nc24722;
wire nc24723;
wire nc24724;
wire nc24725;
wire nc24726;
wire nc24727;
wire nc24728;
wire nc24729;
wire nc24730;
wire nc24731;
wire nc24732;
wire nc24733;
wire nc24734;
wire nc24735;
wire nc24736;
wire nc24737;
wire nc24738;
wire nc24739;
wire nc24740;
wire nc24741;
wire nc24742;
wire nc24743;
wire nc24744;
wire nc24745;
wire nc24746;
wire nc24747;
wire nc24748;
wire nc24749;
wire nc24750;
wire nc24751;
wire nc24752;
wire nc24753;
wire nc24754;
wire nc24755;
wire nc24756;
wire nc24757;
wire nc24758;
wire nc24759;
wire nc24760;
wire nc24761;
wire nc24762;
wire nc24763;
wire nc24764;
wire nc24765;
wire nc24766;
wire nc24767;
wire nc24768;
wire nc24769;
wire nc24770;
wire nc24771;
wire nc24772;
wire nc24773;
wire nc24774;
wire nc24775;
wire nc24776;
wire nc24777;
wire nc24778;
wire nc24779;
wire nc24780;
wire nc24781;
wire nc24782;
wire nc24783;
wire nc24784;
wire nc24785;
wire nc24786;
wire nc24787;
wire nc24788;
wire nc24789;
wire nc24790;
wire nc24791;
wire nc24792;
wire nc24793;
wire nc24794;
wire nc24795;
wire nc24796;
wire nc24797;
wire nc24798;
wire nc24799;
wire nc24800;
wire nc24801;
wire nc24802;
wire nc24803;
wire nc24804;
wire nc24805;
wire nc24806;
wire nc24807;
wire nc24808;
wire nc24809;
wire nc24810;
wire nc24811;
wire nc24812;
wire nc24813;
wire nc24814;
wire nc24815;
wire nc24816;
wire nc24817;
wire nc24818;
wire nc24819;
wire nc24820;
wire nc24821;
wire nc24822;
wire nc24823;
wire nc24824;
wire nc24825;
wire nc24826;
wire nc24827;
wire nc24828;
wire nc24829;
wire nc24830;
wire nc24831;
wire nc24832;
wire nc24833;
wire nc24834;
wire nc24835;
wire nc24836;
wire nc24837;
wire nc24838;
wire nc24839;
wire nc24840;
wire nc24841;
wire nc24842;
wire nc24843;
wire nc24844;
wire nc24845;
wire nc24846;
wire nc24847;
wire nc24848;
wire nc24849;
wire nc24850;
wire nc24851;
wire nc24852;
wire nc24853;
wire nc24854;
wire nc24855;
wire nc24856;
wire nc24857;
wire nc24858;
wire nc24859;
wire nc24860;
wire nc24861;
wire nc24862;
wire nc24863;
wire nc24864;
wire nc24865;
wire nc24866;
wire nc24867;
wire nc24868;
wire nc24869;
wire nc24870;
wire nc24871;
wire nc24872;
wire nc24873;
wire nc24874;
wire nc24875;
wire nc24876;
wire nc24877;
wire nc24878;
wire nc24879;
wire nc24880;
wire nc24881;
wire nc24882;
wire nc24883;
wire nc24884;
wire nc24885;
wire nc24886;
wire nc24887;
wire nc24888;
wire nc24889;
wire nc24890;
wire nc24891;
wire nc24892;
wire nc24893;
wire nc24894;
wire nc24895;
wire nc24896;
wire nc24897;
wire nc24898;
wire nc24899;
wire nc24900;
wire nc24901;
wire nc24902;
wire nc24903;
wire nc24904;
wire nc24905;
wire nc24906;
wire nc24907;
wire nc24908;
wire nc24909;
wire nc24910;
wire nc24911;
wire nc24912;
wire nc24913;
wire nc24914;
wire nc24915;
wire nc24916;
wire nc24917;
wire nc24918;
wire nc24919;
wire nc24920;
wire nc24921;
wire nc24922;
wire nc24923;
wire nc24924;
wire nc24925;
wire nc24926;
wire nc24927;
wire nc24928;
wire nc24929;
wire nc24930;
wire nc24931;
wire nc24932;
wire nc24933;
wire nc24934;
wire nc24935;
wire nc24936;
wire nc24937;
wire nc24938;
wire nc24939;
wire nc24940;
wire nc24941;
wire nc24942;
wire nc24943;
wire nc24944;
wire nc24945;
wire nc24946;
wire nc24947;
wire nc24948;
wire nc24949;
wire nc24950;
wire nc24951;
wire nc24952;
wire nc24953;
wire nc24954;
wire nc24955;
wire nc24956;
wire nc24957;
wire nc24958;
wire nc24959;
wire nc24960;
wire nc24961;
wire nc24962;
wire nc24963;
wire nc24964;
wire nc24965;
wire nc24966;
wire nc24967;
wire nc24968;
wire nc24969;
wire nc24970;
wire nc24971;
wire nc24972;
wire nc24973;
wire nc24974;
wire nc24975;
wire nc24976;
wire nc24977;
wire nc24978;
wire nc24979;
wire nc24980;
wire nc24981;
wire nc24982;
wire nc24983;
wire nc24984;
wire nc24985;
wire nc24986;
wire nc24987;
wire nc24988;
wire nc24989;
wire nc24990;
wire nc24991;
wire nc24992;
wire nc24993;
wire nc24994;
wire nc24995;
wire nc24996;
wire nc24997;
wire nc24998;
wire nc24999;
wire nc25000;
wire nc25001;
wire nc25002;
wire nc25003;
wire nc25004;
wire nc25005;
wire nc25006;
wire nc25007;
wire nc25008;
wire nc25009;
wire nc25010;
wire nc25011;
wire nc25012;
wire nc25013;
wire nc25014;
wire nc25015;
wire nc25016;
wire nc25017;
wire nc25018;
wire nc25019;
wire nc25020;
wire nc25021;
wire nc25022;
wire nc25023;
wire nc25024;
wire nc25025;
wire nc25026;
wire nc25027;
wire nc25028;
wire nc25029;
wire nc25030;
wire nc25031;
wire nc25032;
wire nc25033;
wire nc25034;
wire nc25035;
wire nc25036;
wire nc25037;
wire nc25038;
wire nc25039;
wire nc25040;
wire nc25041;
wire nc25042;
wire nc25043;
wire nc25044;
wire nc25045;
wire nc25046;
wire nc25047;
wire nc25048;
wire nc25049;
wire nc25050;
wire nc25051;
wire nc25052;
wire nc25053;
wire nc25054;
wire nc25055;
wire nc25056;
wire nc25057;
wire nc25058;
wire nc25059;
wire nc25060;
wire nc25061;
wire nc25062;
wire nc25063;
wire nc25064;
wire nc25065;
wire nc25066;
wire nc25067;
wire nc25068;
wire nc25069;
wire nc25070;
wire nc25071;
wire nc25072;
wire nc25073;
wire nc25074;
wire nc25075;
wire nc25076;
wire nc25077;
wire nc25078;
wire nc25079;
wire nc25080;
wire nc25081;
wire nc25082;
wire nc25083;
wire nc25084;
wire nc25085;
wire nc25086;
wire nc25087;
wire nc25088;
wire nc25089;
wire nc25090;
wire nc25091;
wire nc25092;
wire nc25093;
wire nc25094;
wire nc25095;
wire nc25096;
wire nc25097;
wire nc25098;
wire nc25099;
wire nc25100;
wire nc25101;
wire nc25102;
wire nc25103;
wire nc25104;
wire nc25105;
wire nc25106;
wire nc25107;
wire nc25108;
wire nc25109;
wire nc25110;
wire nc25111;
wire nc25112;
wire nc25113;
wire nc25114;
wire nc25115;
wire nc25116;
wire nc25117;
wire nc25118;
wire nc25119;
wire nc25120;
wire nc25121;
wire nc25122;
wire nc25123;
wire nc25124;
wire nc25125;
wire nc25126;
wire nc25127;
wire nc25128;
wire nc25129;
wire nc25130;
wire nc25131;
wire nc25132;
wire nc25133;
wire nc25134;
wire nc25135;
wire nc25136;
wire nc25137;
wire nc25138;
wire nc25139;
wire nc25140;
wire nc25141;
wire nc25142;
wire nc25143;
wire nc25144;
wire nc25145;
wire nc25146;
wire nc25147;
wire nc25148;
wire nc25149;
wire nc25150;
wire nc25151;
wire nc25152;
wire nc25153;
wire nc25154;
wire nc25155;
wire nc25156;
wire nc25157;
wire nc25158;
wire nc25159;
wire nc25160;
wire nc25161;
wire nc25162;
wire nc25163;
wire nc25164;
wire nc25165;
wire nc25166;
wire nc25167;
wire nc25168;
wire nc25169;
wire nc25170;
wire nc25171;
wire nc25172;
wire nc25173;
wire nc25174;
wire nc25175;
wire nc25176;
wire nc25177;
wire nc25178;
wire nc25179;
wire nc25180;
wire nc25181;
wire nc25182;
wire nc25183;
wire nc25184;
wire nc25185;
wire nc25186;
wire nc25187;
wire nc25188;
wire nc25189;
wire nc25190;
wire nc25191;
wire nc25192;
wire nc25193;
wire nc25194;
wire nc25195;
wire nc25196;
wire nc25197;
wire nc25198;
wire nc25199;
wire nc25200;
wire nc25201;
wire nc25202;
wire nc25203;
wire nc25204;
wire nc25205;
wire nc25206;
wire nc25207;
wire nc25208;
wire nc25209;
wire nc25210;
wire nc25211;
wire nc25212;
wire nc25213;
wire nc25214;
wire nc25215;
wire nc25216;
wire nc25217;
wire nc25218;
wire nc25219;
wire nc25220;
wire nc25221;
wire nc25222;
wire nc25223;
wire nc25224;
wire nc25225;
wire nc25226;
wire nc25227;
wire nc25228;
wire nc25229;
wire nc25230;
wire nc25231;
wire nc25232;
wire nc25233;
wire nc25234;
wire nc25235;
wire nc25236;
wire nc25237;
wire nc25238;
wire nc25239;
wire nc25240;
wire nc25241;
wire nc25242;
wire nc25243;
wire nc25244;
wire nc25245;
wire nc25246;
wire nc25247;
wire nc25248;
wire nc25249;
wire nc25250;
wire nc25251;
wire nc25252;
wire nc25253;
wire nc25254;
wire nc25255;
wire nc25256;
wire nc25257;
wire nc25258;
wire nc25259;
wire nc25260;
wire nc25261;
wire nc25262;
wire nc25263;
wire nc25264;
wire nc25265;
wire nc25266;
wire nc25267;
wire nc25268;
wire nc25269;
wire nc25270;
wire nc25271;
wire nc25272;
wire nc25273;
wire nc25274;
wire nc25275;
wire nc25276;
wire nc25277;
wire nc25278;
wire nc25279;
wire nc25280;
wire nc25281;
wire nc25282;
wire nc25283;
wire nc25284;
wire nc25285;
wire nc25286;
wire nc25287;
wire nc25288;
wire nc25289;
wire nc25290;
wire nc25291;
wire nc25292;
wire nc25293;
wire nc25294;
wire nc25295;
wire nc25296;
wire nc25297;
wire nc25298;
wire nc25299;
wire nc25300;
wire nc25301;
wire nc25302;
wire nc25303;
wire nc25304;
wire nc25305;
wire nc25306;
wire nc25307;
wire nc25308;
wire nc25309;
wire nc25310;
wire nc25311;
wire nc25312;
wire nc25313;
wire nc25314;
wire nc25315;
wire nc25316;
wire nc25317;
wire nc25318;
wire nc25319;
wire nc25320;
wire nc25321;
wire nc25322;
wire nc25323;
wire nc25324;
wire nc25325;
wire nc25326;
wire nc25327;
wire nc25328;
wire nc25329;
wire nc25330;
wire nc25331;
wire nc25332;
wire nc25333;
wire nc25334;
wire nc25335;
wire nc25336;
wire nc25337;
wire nc25338;
wire nc25339;
wire nc25340;
wire nc25341;
wire nc25342;
wire nc25343;
wire nc25344;
wire nc25345;
wire nc25346;
wire nc25347;
wire nc25348;
wire nc25349;
wire nc25350;
wire nc25351;
wire nc25352;
wire nc25353;
wire nc25354;
wire nc25355;
wire nc25356;
wire nc25357;
wire nc25358;
wire nc25359;
wire nc25360;
wire nc25361;
wire nc25362;
wire nc25363;
wire nc25364;
wire nc25365;
wire nc25366;
wire nc25367;
wire nc25368;
wire nc25369;
wire nc25370;
wire nc25371;
wire nc25372;
wire nc25373;
wire nc25374;
wire nc25375;
wire nc25376;
wire nc25377;
wire nc25378;
wire nc25379;
wire nc25380;
wire nc25381;
wire nc25382;
wire nc25383;
wire nc25384;
wire nc25385;
wire nc25386;
wire nc25387;
wire nc25388;
wire nc25389;
wire nc25390;
wire nc25391;
wire nc25392;
wire nc25393;
wire nc25394;
wire nc25395;
wire nc25396;
wire nc25397;
wire nc25398;
wire nc25399;
wire nc25400;
wire nc25401;
wire nc25402;
wire nc25403;
wire nc25404;
wire nc25405;
wire nc25406;
wire nc25407;
wire nc25408;
wire nc25409;
wire nc25410;
wire nc25411;
wire nc25412;
wire nc25413;
wire nc25414;
wire nc25415;
wire nc25416;
wire nc25417;
wire nc25418;
wire nc25419;
wire nc25420;
wire nc25421;
wire nc25422;
wire nc25423;
wire nc25424;
wire nc25425;
wire nc25426;
wire nc25427;
wire nc25428;
wire nc25429;
wire nc25430;
wire nc25431;
wire nc25432;
wire nc25433;
wire nc25434;
wire nc25435;
wire nc25436;
wire nc25437;
wire nc25438;
wire nc25439;
wire nc25440;
wire nc25441;
wire nc25442;
wire nc25443;
wire nc25444;
wire nc25445;
wire nc25446;
wire nc25447;
wire nc25448;
wire nc25449;
wire nc25450;
wire nc25451;
wire nc25452;
wire nc25453;
wire nc25454;
wire nc25455;
wire nc25456;
wire nc25457;
wire nc25458;
wire nc25459;
wire nc25460;
wire nc25461;
wire nc25462;
wire nc25463;
wire nc25464;
wire nc25465;
wire nc25466;
wire nc25467;
wire nc25468;
wire nc25469;
wire nc25470;
wire nc25471;
wire nc25472;
wire nc25473;
wire nc25474;
wire nc25475;
wire nc25476;
wire nc25477;
wire nc25478;
wire nc25479;
wire nc25480;
wire nc25481;
wire nc25482;
wire nc25483;
wire nc25484;
wire nc25485;
wire nc25486;
wire nc25487;
wire nc25488;
wire nc25489;
wire nc25490;
wire nc25491;
wire nc25492;
wire nc25493;
wire nc25494;
wire nc25495;
wire nc25496;
wire nc25497;
wire nc25498;
wire nc25499;
wire nc25500;
wire nc25501;
wire nc25502;
wire nc25503;
wire nc25504;
wire nc25505;
wire nc25506;
wire nc25507;
wire nc25508;
wire nc25509;
wire nc25510;
wire nc25511;
wire nc25512;
wire nc25513;
wire nc25514;
wire nc25515;
wire nc25516;
wire nc25517;
wire nc25518;
wire nc25519;
wire nc25520;
wire nc25521;
wire nc25522;
wire nc25523;
wire nc25524;
wire nc25525;
wire nc25526;
wire nc25527;
wire nc25528;
wire nc25529;
wire nc25530;
wire nc25531;
wire nc25532;
wire nc25533;
wire nc25534;
wire nc25535;
wire nc25536;
wire nc25537;
wire nc25538;
wire nc25539;
wire nc25540;
wire nc25541;
wire nc25542;
wire nc25543;
wire nc25544;
wire nc25545;
wire nc25546;
wire nc25547;
wire nc25548;
wire nc25549;
wire nc25550;
wire nc25551;
wire nc25552;
wire nc25553;
wire nc25554;
wire nc25555;
wire nc25556;
wire nc25557;
wire nc25558;
wire nc25559;
wire nc25560;
wire nc25561;
wire nc25562;
wire nc25563;
wire nc25564;
wire nc25565;
wire nc25566;
wire nc25567;
wire nc25568;
wire nc25569;
wire nc25570;
wire nc25571;
wire nc25572;
wire nc25573;
wire nc25574;
wire nc25575;
wire nc25576;
wire nc25577;
wire nc25578;
wire nc25579;
wire nc25580;
wire nc25581;
wire nc25582;
wire nc25583;
wire nc25584;
wire nc25585;
wire nc25586;
wire nc25587;
wire nc25588;
wire nc25589;
wire nc25590;
wire nc25591;
wire nc25592;
wire nc25593;
wire nc25594;
wire nc25595;
wire nc25596;
wire nc25597;
wire nc25598;
wire nc25599;
wire nc25600;
wire nc25601;
wire nc25602;
wire nc25603;
wire nc25604;
wire nc25605;
wire nc25606;
wire nc25607;
wire nc25608;
wire nc25609;
wire nc25610;
wire nc25611;
wire nc25612;
wire nc25613;
wire nc25614;
wire nc25615;
wire nc25616;
wire nc25617;
wire nc25618;
wire nc25619;
wire nc25620;
wire nc25621;
wire nc25622;
wire nc25623;
wire nc25624;
wire nc25625;
wire nc25626;
wire nc25627;
wire nc25628;
wire nc25629;
wire nc25630;
wire nc25631;
wire nc25632;
wire nc25633;
wire nc25634;
wire nc25635;
wire nc25636;
wire nc25637;
wire nc25638;
wire nc25639;
wire nc25640;
wire nc25641;
wire nc25642;
wire nc25643;
wire nc25644;
wire nc25645;
wire nc25646;
wire nc25647;
wire nc25648;
wire nc25649;
wire nc25650;
wire nc25651;
wire nc25652;
wire nc25653;
wire nc25654;
wire nc25655;
wire nc25656;
wire nc25657;
wire nc25658;
wire nc25659;
wire nc25660;
wire nc25661;
wire nc25662;
wire nc25663;
wire nc25664;
wire nc25665;
wire nc25666;
wire nc25667;
wire nc25668;
wire nc25669;
wire nc25670;
wire nc25671;
wire nc25672;
wire nc25673;
wire nc25674;
wire nc25675;
wire nc25676;
wire nc25677;
wire nc25678;
wire nc25679;
wire nc25680;
wire nc25681;
wire nc25682;
wire nc25683;
wire nc25684;
wire nc25685;
wire nc25686;
wire nc25687;
wire nc25688;
wire nc25689;
wire nc25690;
wire nc25691;
wire nc25692;
wire nc25693;
wire nc25694;
wire nc25695;
wire nc25696;
wire nc25697;
wire nc25698;
wire nc25699;
wire nc25700;
wire nc25701;
wire nc25702;
wire nc25703;
wire nc25704;
wire nc25705;
wire nc25706;
wire nc25707;
wire nc25708;
wire nc25709;
wire nc25710;
wire nc25711;
wire nc25712;
wire nc25713;
wire nc25714;
wire nc25715;
wire nc25716;
wire nc25717;
wire nc25718;
wire nc25719;
wire nc25720;
wire nc25721;
wire nc25722;
wire nc25723;
wire nc25724;
wire nc25725;
wire nc25726;
wire nc25727;
wire nc25728;
wire nc25729;
wire nc25730;
wire nc25731;
wire nc25732;
wire nc25733;
wire nc25734;
wire nc25735;
wire nc25736;
wire nc25737;
wire nc25738;
wire nc25739;
wire nc25740;
wire nc25741;
wire nc25742;
wire nc25743;
wire nc25744;
wire nc25745;
wire nc25746;
wire nc25747;
wire nc25748;
wire nc25749;
wire nc25750;
wire nc25751;
wire nc25752;
wire nc25753;
wire nc25754;
wire nc25755;
wire nc25756;
wire nc25757;
wire nc25758;
wire nc25759;
wire nc25760;
wire nc25761;
wire nc25762;
wire nc25763;
wire nc25764;
wire nc25765;
wire nc25766;
wire nc25767;
wire nc25768;
wire nc25769;
wire nc25770;
wire nc25771;
wire nc25772;
wire nc25773;
wire nc25774;
wire nc25775;
wire nc25776;
wire nc25777;
wire nc25778;
wire nc25779;
wire nc25780;
wire nc25781;
wire nc25782;
wire nc25783;
wire nc25784;
wire nc25785;
wire nc25786;
wire nc25787;
wire nc25788;
wire nc25789;
wire nc25790;
wire nc25791;
wire nc25792;
wire nc25793;
wire nc25794;
wire nc25795;
wire nc25796;
wire nc25797;
wire nc25798;
wire nc25799;
wire nc25800;
wire nc25801;
wire nc25802;
wire nc25803;
wire nc25804;
wire nc25805;
wire nc25806;
wire nc25807;
wire nc25808;
wire nc25809;
wire nc25810;
wire nc25811;
wire nc25812;
wire nc25813;
wire nc25814;
wire nc25815;
wire nc25816;
wire nc25817;
wire nc25818;
wire nc25819;
wire nc25820;
wire nc25821;
wire nc25822;
wire nc25823;
wire nc25824;
wire nc25825;
wire nc25826;
wire nc25827;
wire nc25828;
wire nc25829;
wire nc25830;
wire nc25831;
wire nc25832;
wire nc25833;
wire nc25834;
wire nc25835;
wire nc25836;
wire nc25837;
wire nc25838;
wire nc25839;
wire nc25840;
wire nc25841;
wire nc25842;
wire nc25843;
wire nc25844;
wire nc25845;
wire nc25846;
wire nc25847;
wire nc25848;
wire nc25849;
wire nc25850;
wire nc25851;
wire nc25852;
wire nc25853;
wire nc25854;
wire nc25855;
wire nc25856;
wire nc25857;
wire nc25858;
wire nc25859;
wire nc25860;
wire nc25861;
wire nc25862;
wire nc25863;
wire nc25864;
wire nc25865;
wire nc25866;
wire nc25867;
wire nc25868;
wire nc25869;
wire nc25870;
wire nc25871;
wire nc25872;
wire nc25873;
wire nc25874;
wire nc25875;
wire nc25876;
wire nc25877;
wire nc25878;
wire nc25879;
wire nc25880;
wire nc25881;
wire nc25882;
wire nc25883;
wire nc25884;
wire nc25885;
wire nc25886;
wire nc25887;
wire nc25888;
wire nc25889;
wire nc25890;
wire nc25891;
wire nc25892;
wire nc25893;
wire nc25894;
wire nc25895;
wire nc25896;
wire nc25897;
wire nc25898;
wire nc25899;
wire nc25900;
wire nc25901;
wire nc25902;
wire nc25903;
wire nc25904;
wire nc25905;
wire nc25906;
wire nc25907;
wire nc25908;
wire nc25909;
wire nc25910;
wire nc25911;
wire nc25912;
wire nc25913;
wire nc25914;
wire nc25915;
wire nc25916;
wire nc25917;
wire nc25918;
wire nc25919;
wire nc25920;
wire nc25921;
wire nc25922;
wire nc25923;
wire nc25924;
wire nc25925;
wire nc25926;
wire nc25927;
wire nc25928;
wire nc25929;
wire nc25930;
wire nc25931;
wire nc25932;
wire nc25933;
wire nc25934;
wire nc25935;
wire nc25936;
wire nc25937;
wire nc25938;
wire nc25939;
wire nc25940;
wire nc25941;
wire nc25942;
wire nc25943;
wire nc25944;
wire nc25945;
wire nc25946;
wire nc25947;
wire nc25948;
wire nc25949;
wire nc25950;
wire nc25951;
wire nc25952;
wire nc25953;
wire nc25954;
wire nc25955;
wire nc25956;
wire nc25957;
wire nc25958;
wire nc25959;
wire nc25960;
wire nc25961;
wire nc25962;
wire nc25963;
wire nc25964;
wire nc25965;
wire nc25966;
wire nc25967;
wire nc25968;
wire nc25969;
wire nc25970;
wire nc25971;
wire nc25972;
wire nc25973;
wire nc25974;
wire nc25975;
wire nc25976;
wire nc25977;
wire nc25978;
wire nc25979;
wire nc25980;
wire nc25981;
wire nc25982;
wire nc25983;
wire nc25984;
wire nc25985;
wire nc25986;
wire nc25987;
wire nc25988;
wire nc25989;
wire nc25990;
wire nc25991;
wire nc25992;
wire nc25993;
wire nc25994;
wire nc25995;
wire nc25996;
wire nc25997;
wire nc25998;
wire nc25999;
wire nc26000;
wire nc26001;
wire nc26002;
wire nc26003;
wire nc26004;
wire nc26005;
wire nc26006;
wire nc26007;
wire nc26008;
wire nc26009;
wire nc26010;
wire nc26011;
wire nc26012;
wire nc26013;
wire nc26014;
wire nc26015;
wire nc26016;
wire nc26017;
wire nc26018;
wire nc26019;
wire nc26020;
wire nc26021;
wire nc26022;
wire nc26023;
wire nc26024;
wire nc26025;
wire nc26026;
wire nc26027;
wire nc26028;
wire nc26029;
wire nc26030;
wire nc26031;
wire nc26032;
wire nc26033;
wire nc26034;
wire nc26035;
wire nc26036;
wire nc26037;
wire nc26038;
wire nc26039;
wire nc26040;
wire nc26041;
wire nc26042;
wire nc26043;
wire nc26044;
wire nc26045;
wire nc26046;
wire nc26047;
wire nc26048;
wire nc26049;
wire nc26050;
wire nc26051;
wire nc26052;
wire nc26053;
wire nc26054;
wire nc26055;
wire nc26056;
wire nc26057;
wire nc26058;
wire nc26059;
wire nc26060;
wire nc26061;
wire nc26062;
wire nc26063;
wire nc26064;
wire nc26065;
wire nc26066;
wire nc26067;
wire nc26068;
wire nc26069;
wire nc26070;
wire nc26071;
wire nc26072;
wire nc26073;
wire nc26074;
wire nc26075;
wire nc26076;
wire nc26077;
wire nc26078;
wire nc26079;
wire nc26080;
wire nc26081;
wire nc26082;
wire nc26083;
wire nc26084;
wire nc26085;
wire nc26086;
wire nc26087;
wire nc26088;
wire nc26089;
wire nc26090;
wire nc26091;
wire nc26092;
wire nc26093;
wire nc26094;
wire nc26095;
wire nc26096;
wire nc26097;
wire nc26098;
wire nc26099;
wire nc26100;
wire nc26101;
wire nc26102;
wire nc26103;
wire nc26104;
wire nc26105;
wire nc26106;
wire nc26107;
wire nc26108;
wire nc26109;
wire nc26110;
wire nc26111;
wire nc26112;
wire nc26113;
wire nc26114;
wire nc26115;
wire nc26116;
wire nc26117;
wire nc26118;
wire nc26119;
wire nc26120;
wire nc26121;
wire nc26122;
wire nc26123;
wire nc26124;
wire nc26125;
wire nc26126;
wire nc26127;
wire nc26128;
wire nc26129;
wire nc26130;
wire nc26131;
wire nc26132;
wire nc26133;
wire nc26134;
wire nc26135;
wire nc26136;
wire nc26137;
wire nc26138;
wire nc26139;
wire nc26140;
wire nc26141;
wire nc26142;
wire nc26143;
wire nc26144;
wire nc26145;
wire nc26146;
wire nc26147;
wire nc26148;
wire nc26149;
wire nc26150;
wire nc26151;
wire nc26152;
wire nc26153;
wire nc26154;
wire nc26155;
wire nc26156;
wire nc26157;
wire nc26158;
wire nc26159;
wire nc26160;
wire nc26161;
wire nc26162;
wire nc26163;
wire nc26164;
wire nc26165;
wire nc26166;
wire nc26167;
wire nc26168;
wire nc26169;
wire nc26170;
wire nc26171;
wire nc26172;
wire nc26173;
wire nc26174;
wire nc26175;
wire nc26176;
wire nc26177;
wire nc26178;
wire nc26179;
wire nc26180;
wire nc26181;
wire nc26182;
wire nc26183;
wire nc26184;
wire nc26185;
wire nc26186;
wire nc26187;
wire nc26188;
wire nc26189;
wire nc26190;
wire nc26191;
wire nc26192;
wire nc26193;
wire nc26194;
wire nc26195;
wire nc26196;
wire nc26197;
wire nc26198;
wire nc26199;
wire nc26200;
wire nc26201;
wire nc26202;
wire nc26203;
wire nc26204;
wire nc26205;
wire nc26206;
wire nc26207;
wire nc26208;
wire nc26209;
wire nc26210;
wire nc26211;
wire nc26212;
wire nc26213;
wire nc26214;
wire nc26215;
wire nc26216;
wire nc26217;
wire nc26218;
wire nc26219;
wire nc26220;
wire nc26221;
wire nc26222;
wire nc26223;
wire nc26224;
wire nc26225;
wire nc26226;
wire nc26227;
wire nc26228;
wire nc26229;
wire nc26230;
wire nc26231;
wire nc26232;
wire nc26233;
wire nc26234;
wire nc26235;
wire nc26236;
wire nc26237;
wire nc26238;
wire nc26239;
wire nc26240;
wire nc26241;
wire nc26242;
wire nc26243;
wire nc26244;
wire nc26245;
wire nc26246;
wire nc26247;
wire nc26248;
wire nc26249;
wire nc26250;
wire nc26251;
wire nc26252;
wire nc26253;
wire nc26254;
wire nc26255;
wire nc26256;
wire nc26257;
wire nc26258;
wire nc26259;
wire nc26260;
wire nc26261;
wire nc26262;
wire nc26263;
wire nc26264;
wire nc26265;
wire nc26266;
wire nc26267;
wire nc26268;
wire nc26269;
wire nc26270;
wire nc26271;
wire nc26272;
wire nc26273;
wire nc26274;
wire nc26275;
wire nc26276;
wire nc26277;
wire nc26278;
wire nc26279;
wire nc26280;
wire nc26281;
wire nc26282;
wire nc26283;
wire nc26284;
wire nc26285;
wire nc26286;
wire nc26287;
wire nc26288;
wire nc26289;
wire nc26290;
wire nc26291;
wire nc26292;
wire nc26293;
wire nc26294;
wire nc26295;
wire nc26296;
wire nc26297;
wire nc26298;
wire nc26299;
wire nc26300;
wire nc26301;
wire nc26302;
wire nc26303;
wire nc26304;
wire nc26305;
wire nc26306;
wire nc26307;
wire nc26308;
wire nc26309;
wire nc26310;
wire nc26311;
wire nc26312;
wire nc26313;
wire nc26314;
wire nc26315;
wire nc26316;
wire nc26317;
wire nc26318;
wire nc26319;
wire nc26320;
wire nc26321;
wire nc26322;
wire nc26323;
wire nc26324;
wire nc26325;
wire nc26326;
wire nc26327;
wire nc26328;
wire nc26329;
wire nc26330;
wire nc26331;
wire nc26332;
wire nc26333;
wire nc26334;
wire nc26335;
wire nc26336;
wire nc26337;
wire nc26338;
wire nc26339;
wire nc26340;
wire nc26341;
wire nc26342;
wire nc26343;
wire nc26344;
wire nc26345;
wire nc26346;
wire nc26347;
wire nc26348;
wire nc26349;
wire nc26350;
wire nc26351;
wire nc26352;
wire nc26353;
wire nc26354;
wire nc26355;
wire nc26356;
wire nc26357;
wire nc26358;
wire nc26359;
wire nc26360;
wire nc26361;
wire nc26362;
wire nc26363;
wire nc26364;
wire nc26365;
wire nc26366;
wire nc26367;
wire nc26368;
wire nc26369;
wire nc26370;
wire nc26371;
wire nc26372;
wire nc26373;
wire nc26374;
wire nc26375;
wire nc26376;
wire nc26377;
wire nc26378;
wire nc26379;
wire nc26380;
wire nc26381;
wire nc26382;
wire nc26383;
wire nc26384;
wire nc26385;
wire nc26386;
wire nc26387;
wire nc26388;
wire nc26389;
wire nc26390;
wire nc26391;
wire nc26392;
wire nc26393;
wire nc26394;
wire nc26395;
wire nc26396;
wire nc26397;
wire nc26398;
wire nc26399;
wire nc26400;
wire nc26401;
wire nc26402;
wire nc26403;
wire nc26404;
wire nc26405;
wire nc26406;
wire nc26407;
wire nc26408;
wire nc26409;
wire nc26410;
wire nc26411;
wire nc26412;
wire nc26413;
wire nc26414;
wire nc26415;
wire nc26416;
wire nc26417;
wire nc26418;
wire nc26419;
wire nc26420;
wire nc26421;
wire nc26422;
wire nc26423;
wire nc26424;
wire nc26425;
wire nc26426;
wire nc26427;
wire nc26428;
wire nc26429;
wire nc26430;
wire nc26431;
wire nc26432;
wire nc26433;
wire nc26434;
wire nc26435;
wire nc26436;
wire nc26437;
wire nc26438;
wire nc26439;
wire nc26440;
wire nc26441;
wire nc26442;
wire nc26443;
wire nc26444;
wire nc26445;
wire nc26446;
wire nc26447;
wire nc26448;
wire nc26449;
wire nc26450;
wire nc26451;
wire nc26452;
wire nc26453;
wire nc26454;
wire nc26455;
wire nc26456;
wire nc26457;
wire nc26458;
wire nc26459;
wire nc26460;
wire nc26461;
wire nc26462;
wire nc26463;
wire nc26464;
wire nc26465;
wire nc26466;
wire nc26467;
wire nc26468;
wire nc26469;
wire nc26470;
wire nc26471;
wire nc26472;
wire nc26473;
wire nc26474;
wire nc26475;
wire nc26476;
wire nc26477;
wire nc26478;
wire nc26479;
wire nc26480;
wire nc26481;
wire nc26482;
wire nc26483;
wire nc26484;
wire nc26485;
wire nc26486;
wire nc26487;
wire nc26488;
wire nc26489;
wire nc26490;
wire nc26491;
wire nc26492;
wire nc26493;
wire nc26494;
wire nc26495;
wire nc26496;
wire nc26497;
wire nc26498;
wire nc26499;
wire nc26500;
wire nc26501;
wire nc26502;
wire nc26503;
wire nc26504;
wire nc26505;
wire nc26506;
wire nc26507;
wire nc26508;
wire nc26509;
wire nc26510;
wire nc26511;
wire nc26512;
wire nc26513;
wire nc26514;
wire nc26515;
wire nc26516;
wire nc26517;
wire nc26518;
wire nc26519;
wire nc26520;
wire nc26521;
wire nc26522;
wire nc26523;
wire nc26524;
wire nc26525;
wire nc26526;
wire nc26527;
wire nc26528;
wire nc26529;
wire nc26530;
wire nc26531;
wire nc26532;
wire nc26533;
wire nc26534;
wire nc26535;
wire nc26536;
wire nc26537;
wire nc26538;
wire nc26539;
wire nc26540;
wire nc26541;
wire nc26542;
wire nc26543;
wire nc26544;
wire nc26545;
wire nc26546;
wire nc26547;
wire nc26548;
wire nc26549;
wire nc26550;
wire nc26551;
wire nc26552;
wire nc26553;
wire nc26554;
wire nc26555;
wire nc26556;
wire nc26557;
wire nc26558;
wire nc26559;
wire nc26560;
wire nc26561;
wire nc26562;
wire nc26563;
wire nc26564;
wire nc26565;
wire nc26566;
wire nc26567;
wire nc26568;
wire nc26569;
wire nc26570;
wire nc26571;
wire nc26572;
wire nc26573;
wire nc26574;
wire nc26575;
wire nc26576;
wire nc26577;
wire nc26578;
wire nc26579;
wire nc26580;
wire nc26581;
wire nc26582;
wire nc26583;
wire nc26584;
wire nc26585;
wire nc26586;
wire nc26587;
wire nc26588;
wire nc26589;
wire nc26590;
wire nc26591;
wire nc26592;
wire nc26593;
wire nc26594;
wire nc26595;
wire nc26596;
wire nc26597;
wire nc26598;
wire nc26599;
wire nc26600;
wire nc26601;
wire nc26602;
wire nc26603;
wire nc26604;
wire nc26605;
wire nc26606;
wire nc26607;
wire nc26608;
wire nc26609;
wire nc26610;
wire nc26611;
wire nc26612;
wire nc26613;
wire nc26614;
wire nc26615;
wire nc26616;
wire nc26617;
wire nc26618;
wire nc26619;
wire nc26620;
wire nc26621;
wire nc26622;
wire nc26623;
wire nc26624;
wire nc26625;
wire nc26626;
wire nc26627;
wire nc26628;
wire nc26629;
wire nc26630;
wire nc26631;
wire nc26632;
wire nc26633;
wire nc26634;
wire nc26635;
wire nc26636;
wire nc26637;
wire nc26638;
wire nc26639;
wire nc26640;
wire nc26641;
wire nc26642;
wire nc26643;
wire nc26644;
wire nc26645;
wire nc26646;
wire nc26647;
wire nc26648;
wire nc26649;
wire nc26650;
wire nc26651;
wire nc26652;
wire nc26653;
wire nc26654;
wire nc26655;
wire nc26656;
wire nc26657;
wire nc26658;
wire nc26659;
wire nc26660;
wire nc26661;
wire nc26662;
wire nc26663;
wire nc26664;
wire nc26665;
wire nc26666;
wire nc26667;
wire nc26668;
wire nc26669;
wire nc26670;
wire nc26671;
wire nc26672;
wire nc26673;
wire nc26674;
wire nc26675;
wire nc26676;
wire nc26677;
wire nc26678;
wire nc26679;
wire nc26680;
wire nc26681;
wire nc26682;
wire nc26683;
wire nc26684;
wire nc26685;
wire nc26686;
wire nc26687;
wire nc26688;
wire nc26689;
wire nc26690;
wire nc26691;
wire nc26692;
wire nc26693;
wire nc26694;
wire nc26695;
wire nc26696;
wire nc26697;
wire nc26698;
wire nc26699;
wire nc26700;
wire nc26701;
wire nc26702;
wire nc26703;
wire nc26704;
wire nc26705;
wire nc26706;
wire nc26707;
wire nc26708;
wire nc26709;
wire nc26710;
wire nc26711;
wire nc26712;
wire nc26713;
wire nc26714;
wire nc26715;
wire nc26716;
wire nc26717;
wire nc26718;
wire nc26719;
wire nc26720;
wire nc26721;
wire nc26722;
wire nc26723;
wire nc26724;
wire nc26725;
wire nc26726;
wire nc26727;
wire nc26728;
wire nc26729;
wire nc26730;
wire nc26731;
wire nc26732;
wire nc26733;
wire nc26734;
wire nc26735;
wire nc26736;
wire nc26737;
wire nc26738;
wire nc26739;
wire nc26740;
wire nc26741;
wire nc26742;
wire nc26743;
wire nc26744;
wire nc26745;
wire nc26746;
wire nc26747;
wire nc26748;
wire nc26749;
wire nc26750;
wire nc26751;
wire nc26752;
wire nc26753;
wire nc26754;
wire nc26755;
wire nc26756;
wire nc26757;
wire nc26758;
wire nc26759;
wire nc26760;
wire nc26761;
wire nc26762;
wire nc26763;
wire nc26764;
wire nc26765;
wire nc26766;
wire nc26767;
wire nc26768;
wire nc26769;
wire nc26770;
wire nc26771;
wire nc26772;
wire nc26773;
wire nc26774;
wire nc26775;
wire nc26776;
wire nc26777;
wire nc26778;
wire nc26779;
wire nc26780;
wire nc26781;
wire nc26782;
wire nc26783;
wire nc26784;
wire nc26785;
wire nc26786;
wire nc26787;
wire nc26788;
wire nc26789;
wire nc26790;
wire nc26791;
wire nc26792;
wire nc26793;
wire nc26794;
wire nc26795;
wire nc26796;
wire nc26797;
wire nc26798;
wire nc26799;
wire nc26800;
wire nc26801;
wire nc26802;
wire nc26803;
wire nc26804;
wire nc26805;
wire nc26806;
wire nc26807;
wire nc26808;
wire nc26809;
wire nc26810;
wire nc26811;
wire nc26812;
wire nc26813;
wire nc26814;
wire nc26815;
wire nc26816;
wire nc26817;
wire nc26818;
wire nc26819;
wire nc26820;
wire nc26821;
wire nc26822;
wire nc26823;
wire nc26824;
wire nc26825;
wire nc26826;
wire nc26827;
wire nc26828;
wire nc26829;
wire nc26830;
wire nc26831;
wire nc26832;
wire nc26833;
wire nc26834;
wire nc26835;
wire nc26836;
wire nc26837;
wire nc26838;
wire nc26839;
wire nc26840;
wire nc26841;
wire nc26842;
wire nc26843;
wire nc26844;
wire nc26845;
wire nc26846;
wire nc26847;
wire nc26848;
wire nc26849;
wire nc26850;
wire nc26851;
wire nc26852;
wire nc26853;
wire nc26854;
wire nc26855;
wire nc26856;
wire nc26857;
wire nc26858;
wire nc26859;
wire nc26860;
wire nc26861;
wire nc26862;
wire nc26863;
wire nc26864;
wire nc26865;
wire nc26866;
wire nc26867;
wire nc26868;
wire nc26869;
wire nc26870;
wire nc26871;
wire nc26872;
wire nc26873;
wire nc26874;
wire nc26875;
wire nc26876;
wire nc26877;
wire nc26878;
wire nc26879;
wire nc26880;
wire nc26881;
wire nc26882;
wire nc26883;
wire nc26884;
wire nc26885;
wire nc26886;
wire nc26887;
wire nc26888;
wire nc26889;
wire nc26890;
wire nc26891;
wire nc26892;
wire nc26893;
wire nc26894;
wire nc26895;
wire nc26896;
wire nc26897;
wire nc26898;
wire nc26899;
wire nc26900;
wire nc26901;
wire nc26902;
wire nc26903;
wire nc26904;
wire nc26905;
wire nc26906;
wire nc26907;
wire nc26908;
wire nc26909;
wire nc26910;
wire nc26911;
wire nc26912;
wire nc26913;
wire nc26914;
wire nc26915;
wire nc26916;
wire nc26917;
wire nc26918;
wire nc26919;
wire nc26920;
wire nc26921;
wire nc26922;
wire nc26923;
wire nc26924;
wire nc26925;
wire nc26926;
wire nc26927;
wire nc26928;
wire nc26929;
wire nc26930;
wire nc26931;
wire nc26932;
wire nc26933;
wire nc26934;
wire nc26935;
wire nc26936;
wire nc26937;
wire nc26938;
wire nc26939;
wire nc26940;
wire nc26941;
wire nc26942;
wire nc26943;
wire nc26944;
wire nc26945;
wire nc26946;
wire nc26947;
wire nc26948;
wire nc26949;
wire nc26950;
wire nc26951;
wire nc26952;
wire nc26953;
wire nc26954;
wire nc26955;
wire nc26956;
wire nc26957;
wire nc26958;
wire nc26959;
wire nc26960;
wire nc26961;
wire nc26962;
wire nc26963;
wire nc26964;
wire nc26965;
wire nc26966;
wire nc26967;
wire nc26968;
wire nc26969;
wire nc26970;
wire nc26971;
wire nc26972;
wire nc26973;
wire nc26974;
wire nc26975;
wire nc26976;
wire nc26977;
wire nc26978;
wire nc26979;
wire nc26980;
wire nc26981;
wire nc26982;
wire nc26983;
wire nc26984;
wire nc26985;
wire nc26986;
wire nc26987;
wire nc26988;
wire nc26989;
wire nc26990;
wire nc26991;
wire nc26992;
wire nc26993;
wire nc26994;
wire nc26995;
wire nc26996;
wire nc26997;
wire nc26998;
wire nc26999;
wire nc27000;
wire nc27001;
wire nc27002;
wire nc27003;
wire nc27004;
wire nc27005;
wire nc27006;
wire nc27007;
wire nc27008;
wire nc27009;
wire nc27010;
wire nc27011;
wire nc27012;
wire nc27013;
wire nc27014;
wire nc27015;
wire nc27016;
wire nc27017;
wire nc27018;
wire nc27019;
wire nc27020;
wire nc27021;
wire nc27022;
wire nc27023;
wire nc27024;
wire nc27025;
wire nc27026;
wire nc27027;
wire nc27028;
wire nc27029;
wire nc27030;
wire nc27031;
wire nc27032;
wire nc27033;
wire nc27034;
wire nc27035;
wire nc27036;
wire nc27037;
wire nc27038;
wire nc27039;
wire nc27040;
wire nc27041;
wire nc27042;
wire nc27043;
wire nc27044;
wire nc27045;
wire nc27046;
wire nc27047;
wire nc27048;
wire nc27049;
wire nc27050;
wire nc27051;
wire nc27052;
wire nc27053;
wire nc27054;
wire nc27055;
wire nc27056;
wire nc27057;
wire nc27058;
wire nc27059;
wire nc27060;
wire nc27061;
wire nc27062;
wire nc27063;
wire nc27064;
wire nc27065;
wire nc27066;
wire nc27067;
wire nc27068;
wire nc27069;
wire nc27070;
wire nc27071;
wire nc27072;
wire nc27073;
wire nc27074;
wire nc27075;
wire nc27076;
wire nc27077;
wire nc27078;
wire nc27079;
wire nc27080;
wire nc27081;
wire nc27082;
wire nc27083;
wire nc27084;
wire nc27085;
wire nc27086;
wire nc27087;
wire nc27088;
wire nc27089;
wire nc27090;
wire nc27091;
wire nc27092;
wire nc27093;
wire nc27094;
wire nc27095;
wire nc27096;
wire nc27097;
wire nc27098;
wire nc27099;
wire nc27100;
wire nc27101;
wire nc27102;
wire nc27103;
wire nc27104;
wire nc27105;
wire nc27106;
wire nc27107;
wire nc27108;
wire nc27109;
wire nc27110;
wire nc27111;
wire nc27112;
wire nc27113;
wire nc27114;
wire nc27115;
wire nc27116;
wire nc27117;
wire nc27118;
wire nc27119;
wire nc27120;
wire nc27121;
wire nc27122;
wire nc27123;
wire nc27124;
wire nc27125;
wire nc27126;
wire nc27127;
wire nc27128;
wire nc27129;
wire nc27130;
wire nc27131;
wire nc27132;
wire nc27133;
wire nc27134;
wire nc27135;
wire nc27136;
wire nc27137;
wire nc27138;
wire nc27139;
wire nc27140;
wire nc27141;
wire nc27142;
wire nc27143;
wire nc27144;
wire nc27145;
wire nc27146;
wire nc27147;
wire nc27148;
wire nc27149;
wire nc27150;
wire nc27151;
wire nc27152;
wire nc27153;
wire nc27154;
wire nc27155;
wire nc27156;
wire nc27157;
wire nc27158;
wire nc27159;
wire nc27160;
wire nc27161;
wire nc27162;
wire nc27163;
wire nc27164;
wire nc27165;
wire nc27166;
wire nc27167;
wire nc27168;
wire nc27169;
wire nc27170;
wire nc27171;
wire nc27172;
wire nc27173;
wire nc27174;
wire nc27175;
wire nc27176;
wire nc27177;
wire nc27178;
wire nc27179;
wire nc27180;
wire nc27181;
wire nc27182;
wire nc27183;
wire nc27184;
wire nc27185;
wire nc27186;
wire nc27187;
wire nc27188;
wire nc27189;
wire nc27190;
wire nc27191;
wire nc27192;
wire nc27193;
wire nc27194;
wire nc27195;
wire nc27196;
wire nc27197;
wire nc27198;
wire nc27199;
wire nc27200;
wire nc27201;
wire nc27202;
wire nc27203;
wire nc27204;
wire nc27205;
wire nc27206;
wire nc27207;
wire nc27208;
wire nc27209;
wire nc27210;
wire nc27211;
wire nc27212;
wire nc27213;
wire nc27214;
wire nc27215;
wire nc27216;
wire nc27217;
wire nc27218;
wire nc27219;
wire nc27220;
wire nc27221;
wire nc27222;
wire nc27223;
wire nc27224;
wire nc27225;
wire nc27226;
wire nc27227;
wire nc27228;
wire nc27229;
wire nc27230;
wire nc27231;
wire nc27232;
wire nc27233;
wire nc27234;
wire nc27235;
wire nc27236;
wire nc27237;
wire nc27238;
wire nc27239;
wire nc27240;
wire nc27241;
wire nc27242;
wire nc27243;
wire nc27244;
wire nc27245;
wire nc27246;
wire nc27247;
wire nc27248;
wire nc27249;
wire nc27250;
wire nc27251;
wire nc27252;
wire nc27253;
wire nc27254;
wire nc27255;
wire nc27256;
wire nc27257;
wire nc27258;
wire nc27259;
wire nc27260;
wire nc27261;
wire nc27262;
wire nc27263;
wire nc27264;
wire nc27265;
wire nc27266;
wire nc27267;
wire nc27268;
wire nc27269;
wire nc27270;
wire nc27271;
wire nc27272;
wire nc27273;
wire nc27274;
wire nc27275;
wire nc27276;
wire nc27277;
wire nc27278;
wire nc27279;
wire nc27280;
wire nc27281;
wire nc27282;
wire nc27283;
wire nc27284;
wire nc27285;
wire nc27286;
wire nc27287;
wire nc27288;
wire nc27289;
wire nc27290;
wire nc27291;
wire nc27292;
wire nc27293;
wire nc27294;
wire nc27295;
wire nc27296;
wire nc27297;
wire nc27298;
wire nc27299;
wire nc27300;
wire nc27301;
wire nc27302;
wire nc27303;
wire nc27304;
wire nc27305;
wire nc27306;
wire nc27307;
wire nc27308;
wire nc27309;
wire nc27310;
wire nc27311;
wire nc27312;
wire nc27313;
wire nc27314;
wire nc27315;
wire nc27316;
wire nc27317;
wire nc27318;
wire nc27319;
wire nc27320;
wire nc27321;
wire nc27322;
wire nc27323;
wire nc27324;
wire nc27325;
wire nc27326;
wire nc27327;
wire nc27328;
wire nc27329;
wire nc27330;
wire nc27331;
wire nc27332;
wire nc27333;
wire nc27334;
wire nc27335;
wire nc27336;
wire nc27337;
wire nc27338;
wire nc27339;
wire nc27340;
wire nc27341;
wire nc27342;
wire nc27343;
wire nc27344;
wire nc27345;
wire nc27346;
wire nc27347;
wire nc27348;
wire nc27349;
wire nc27350;
wire nc27351;
wire nc27352;
wire nc27353;
wire nc27354;
wire nc27355;
wire nc27356;
wire nc27357;
wire nc27358;
wire nc27359;
wire nc27360;
wire nc27361;
wire nc27362;
wire nc27363;
wire nc27364;
wire nc27365;
wire nc27366;
wire nc27367;
wire nc27368;
wire nc27369;
wire nc27370;
wire nc27371;
wire nc27372;
wire nc27373;
wire nc27374;
wire nc27375;
wire nc27376;
wire nc27377;
wire nc27378;
wire nc27379;
wire nc27380;
wire nc27381;
wire nc27382;
wire nc27383;
wire nc27384;
wire nc27385;
wire nc27386;
wire nc27387;
wire nc27388;
wire nc27389;
wire nc27390;
wire nc27391;
wire nc27392;
wire nc27393;
wire nc27394;
wire nc27395;
wire nc27396;
wire nc27397;
wire nc27398;
wire nc27399;
wire nc27400;
wire nc27401;
wire nc27402;
wire nc27403;
wire nc27404;
wire nc27405;
wire nc27406;
wire nc27407;
wire nc27408;
wire nc27409;
wire nc27410;
wire nc27411;
wire nc27412;
wire nc27413;
wire nc27414;
wire nc27415;
wire nc27416;
wire nc27417;
wire nc27418;
wire nc27419;
wire nc27420;
wire nc27421;
wire nc27422;
wire nc27423;
wire nc27424;
wire nc27425;
wire nc27426;
wire nc27427;
wire nc27428;
wire nc27429;
wire nc27430;
wire nc27431;
wire nc27432;
wire nc27433;
wire nc27434;
wire nc27435;
wire nc27436;
wire nc27437;
wire nc27438;
wire nc27439;
wire nc27440;
wire nc27441;
wire nc27442;
wire nc27443;
wire nc27444;
wire nc27445;
wire nc27446;
wire nc27447;
wire nc27448;
wire nc27449;
wire nc27450;
wire nc27451;
wire nc27452;
wire nc27453;
wire nc27454;
wire nc27455;
wire nc27456;
wire nc27457;
wire nc27458;
wire nc27459;
wire nc27460;
wire nc27461;
wire nc27462;
wire nc27463;
wire nc27464;
wire nc27465;
wire nc27466;
wire nc27467;
wire nc27468;
wire nc27469;
wire nc27470;
wire nc27471;
wire nc27472;
wire nc27473;
wire nc27474;
wire nc27475;
wire nc27476;
wire nc27477;
wire nc27478;
wire nc27479;
wire nc27480;
wire nc27481;
wire nc27482;
wire nc27483;
wire nc27484;
wire nc27485;
wire nc27486;
wire nc27487;
wire nc27488;
wire nc27489;
wire nc27490;
wire nc27491;
wire nc27492;
wire nc27493;
wire nc27494;
wire nc27495;
wire nc27496;
wire nc27497;
wire nc27498;
wire nc27499;
wire nc27500;
wire nc27501;
wire nc27502;
wire nc27503;
wire nc27504;
wire nc27505;
wire nc27506;
wire nc27507;
wire nc27508;
wire nc27509;
wire nc27510;
wire nc27511;
wire nc27512;
wire nc27513;
wire nc27514;
wire nc27515;
wire nc27516;
wire nc27517;
wire nc27518;
wire nc27519;
wire nc27520;
wire nc27521;
wire nc27522;
wire nc27523;
wire nc27524;
wire nc27525;
wire nc27526;
wire nc27527;
wire nc27528;
wire nc27529;
wire nc27530;
wire nc27531;
wire nc27532;
wire nc27533;
wire nc27534;
wire nc27535;
wire nc27536;
wire nc27537;
wire nc27538;
wire nc27539;
wire nc27540;
wire nc27541;
wire nc27542;
wire nc27543;
wire nc27544;
wire nc27545;
wire nc27546;
wire nc27547;
wire nc27548;
wire nc27549;
wire nc27550;
wire nc27551;
wire nc27552;
wire nc27553;
wire nc27554;
wire nc27555;
wire nc27556;
wire nc27557;
wire nc27558;
wire nc27559;
wire nc27560;
wire nc27561;
wire nc27562;
wire nc27563;
wire nc27564;
wire nc27565;
wire nc27566;
wire nc27567;
wire nc27568;
wire nc27569;
wire nc27570;
wire nc27571;
wire nc27572;
wire nc27573;
wire nc27574;
wire nc27575;
wire nc27576;
wire nc27577;
wire nc27578;
wire nc27579;
wire nc27580;
wire nc27581;
wire nc27582;
wire nc27583;
wire nc27584;
wire nc27585;
wire nc27586;
wire nc27587;
wire nc27588;
wire nc27589;
wire nc27590;
wire nc27591;
wire nc27592;
wire nc27593;
wire nc27594;
wire nc27595;
wire nc27596;
wire nc27597;
wire nc27598;
wire nc27599;
wire nc27600;
wire nc27601;
wire nc27602;
wire nc27603;
wire nc27604;
wire nc27605;
wire nc27606;
wire nc27607;
wire nc27608;
wire nc27609;
wire nc27610;
wire nc27611;
wire nc27612;
wire nc27613;
wire nc27614;
wire nc27615;
wire nc27616;
wire nc27617;
wire nc27618;
wire nc27619;
wire nc27620;
wire nc27621;
wire nc27622;
wire nc27623;
wire nc27624;
wire nc27625;
wire nc27626;
wire nc27627;
wire nc27628;
wire nc27629;
wire nc27630;
wire nc27631;
wire nc27632;
wire nc27633;
wire nc27634;
wire nc27635;
wire nc27636;
wire nc27637;
wire nc27638;
wire nc27639;
wire nc27640;
wire nc27641;
wire nc27642;
wire nc27643;
wire nc27644;
wire nc27645;
wire nc27646;
wire nc27647;
wire nc27648;
wire nc27649;
wire nc27650;
wire nc27651;
wire nc27652;
wire nc27653;
wire nc27654;
wire nc27655;
wire nc27656;
wire nc27657;
wire nc27658;
wire nc27659;
wire nc27660;
wire nc27661;
wire nc27662;
wire nc27663;
wire nc27664;
wire nc27665;
wire nc27666;
wire nc27667;
wire nc27668;
wire nc27669;
wire nc27670;
wire nc27671;
wire nc27672;
wire nc27673;
wire nc27674;
wire nc27675;
wire nc27676;
wire nc27677;
wire nc27678;
wire nc27679;
wire nc27680;
wire nc27681;
wire nc27682;
wire nc27683;
wire nc27684;
wire nc27685;
wire nc27686;
wire nc27687;
wire nc27688;
wire nc27689;
wire nc27690;
wire nc27691;
wire nc27692;
wire nc27693;
wire nc27694;
wire nc27695;
wire nc27696;
wire nc27697;
wire nc27698;
wire nc27699;
wire nc27700;
wire nc27701;
wire nc27702;
wire nc27703;
wire nc27704;
wire nc27705;
wire nc27706;
wire nc27707;
wire nc27708;
wire nc27709;
wire nc27710;
wire nc27711;
wire nc27712;
wire nc27713;
wire nc27714;
wire nc27715;
wire nc27716;
wire nc27717;
wire nc27718;
wire nc27719;
wire nc27720;
wire nc27721;
wire nc27722;
wire nc27723;
wire nc27724;
wire nc27725;
wire nc27726;
wire nc27727;
wire nc27728;
wire nc27729;
wire nc27730;
wire nc27731;
wire nc27732;
wire nc27733;
wire nc27734;
wire nc27735;
wire nc27736;
wire nc27737;
wire nc27738;
wire nc27739;
wire nc27740;
wire nc27741;
wire nc27742;
wire nc27743;
wire nc27744;
wire nc27745;
wire nc27746;
wire nc27747;
wire nc27748;
wire nc27749;
wire nc27750;
wire nc27751;
wire nc27752;
wire nc27753;
wire nc27754;
wire nc27755;
wire nc27756;
wire nc27757;
wire nc27758;
wire nc27759;
wire nc27760;
wire nc27761;
wire nc27762;
wire nc27763;
wire nc27764;
wire nc27765;
wire nc27766;
wire nc27767;
wire nc27768;
wire nc27769;
wire nc27770;
wire nc27771;
wire nc27772;
wire nc27773;
wire nc27774;
wire nc27775;
wire nc27776;
wire nc27777;
wire nc27778;
wire nc27779;
wire nc27780;
wire nc27781;
wire nc27782;
wire nc27783;
wire nc27784;
wire nc27785;
wire nc27786;
wire nc27787;
wire nc27788;
wire nc27789;
wire nc27790;
wire nc27791;
wire nc27792;
wire nc27793;
wire nc27794;
wire nc27795;
wire nc27796;
wire nc27797;
wire nc27798;
wire nc27799;
wire nc27800;
wire nc27801;
wire nc27802;
wire nc27803;
wire nc27804;
wire nc27805;
wire nc27806;
wire nc27807;
wire nc27808;
wire nc27809;
wire nc27810;
wire nc27811;
wire nc27812;
wire nc27813;
wire nc27814;
wire nc27815;
wire nc27816;
wire nc27817;
wire nc27818;
wire nc27819;
wire nc27820;
wire nc27821;
wire nc27822;
wire nc27823;
wire nc27824;
wire nc27825;
wire nc27826;
wire nc27827;
wire nc27828;
wire nc27829;
wire nc27830;
wire nc27831;
wire nc27832;
wire nc27833;
wire nc27834;
wire nc27835;
wire nc27836;
wire nc27837;
wire nc27838;
wire nc27839;
wire nc27840;
wire nc27841;
wire nc27842;
wire nc27843;
wire nc27844;
wire nc27845;
wire nc27846;
wire nc27847;
wire nc27848;
wire nc27849;
wire nc27850;
wire nc27851;
wire nc27852;
wire nc27853;
wire nc27854;
wire nc27855;
wire nc27856;
wire nc27857;
wire nc27858;
wire nc27859;
wire nc27860;
wire nc27861;
wire nc27862;
wire nc27863;
wire nc27864;
wire nc27865;
wire nc27866;
wire nc27867;
wire nc27868;
wire nc27869;
wire nc27870;
wire nc27871;
wire nc27872;
wire nc27873;
wire nc27874;
wire nc27875;
wire nc27876;
wire nc27877;
wire nc27878;
wire nc27879;
wire nc27880;
wire nc27881;
wire nc27882;
wire nc27883;
wire nc27884;
wire nc27885;
wire nc27886;
wire nc27887;
wire nc27888;
wire nc27889;
wire nc27890;
wire nc27891;
wire nc27892;
wire nc27893;
wire nc27894;
wire nc27895;
wire nc27896;
wire nc27897;
wire nc27898;
wire nc27899;
wire nc27900;
wire nc27901;
wire nc27902;
wire nc27903;
wire nc27904;
wire nc27905;
wire nc27906;
wire nc27907;
wire nc27908;
wire nc27909;
wire nc27910;
wire nc27911;
wire nc27912;
wire nc27913;
wire nc27914;
wire nc27915;
wire nc27916;
wire nc27917;
wire nc27918;
wire nc27919;
wire nc27920;
wire nc27921;
wire nc27922;
wire nc27923;
wire nc27924;
wire nc27925;
wire nc27926;
wire nc27927;
wire nc27928;
wire nc27929;
wire nc27930;
wire nc27931;
wire nc27932;
wire nc27933;
wire nc27934;
wire nc27935;
wire nc27936;
wire nc27937;
wire nc27938;
wire nc27939;
wire nc27940;
wire nc27941;
wire nc27942;
wire nc27943;
wire nc27944;
wire nc27945;
wire nc27946;
wire nc27947;
wire nc27948;
wire nc27949;
wire nc27950;
wire nc27951;
wire nc27952;
wire nc27953;
wire nc27954;
wire nc27955;
wire nc27956;
wire nc27957;
wire nc27958;
wire nc27959;
wire nc27960;
wire nc27961;
wire nc27962;
wire nc27963;
wire nc27964;
wire nc27965;
wire nc27966;
wire nc27967;
wire nc27968;
wire nc27969;
wire nc27970;
wire nc27971;
wire nc27972;
wire nc27973;
wire nc27974;
wire nc27975;
wire nc27976;
wire nc27977;
wire nc27978;
wire nc27979;
wire nc27980;
wire nc27981;
wire nc27982;
wire nc27983;
wire nc27984;
wire nc27985;
wire nc27986;
wire nc27987;
wire nc27988;
wire nc27989;
wire nc27990;
wire nc27991;
wire nc27992;
wire nc27993;
wire nc27994;
wire nc27995;
wire nc27996;
wire nc27997;
wire nc27998;
wire nc27999;
wire nc28000;
wire nc28001;
wire nc28002;
wire nc28003;
wire nc28004;
wire nc28005;
wire nc28006;
wire nc28007;
wire nc28008;
wire nc28009;
wire nc28010;
wire nc28011;
wire nc28012;
wire nc28013;
wire nc28014;
wire nc28015;
wire nc28016;
wire nc28017;
wire nc28018;
wire nc28019;
wire nc28020;
wire nc28021;
wire nc28022;
wire nc28023;
wire nc28024;
wire nc28025;
wire nc28026;
wire nc28027;
wire nc28028;
wire nc28029;
wire nc28030;
wire nc28031;
wire nc28032;
wire nc28033;
wire nc28034;
wire nc28035;
wire nc28036;
wire nc28037;
wire nc28038;
wire nc28039;
wire nc28040;
wire nc28041;
wire nc28042;
wire nc28043;
wire nc28044;
wire nc28045;
wire nc28046;
wire nc28047;
wire nc28048;
wire nc28049;
wire nc28050;
wire nc28051;
wire nc28052;
wire nc28053;
wire nc28054;
wire nc28055;
wire nc28056;
wire nc28057;
wire nc28058;
wire nc28059;
wire nc28060;
wire nc28061;
wire nc28062;
wire nc28063;
wire nc28064;
wire nc28065;
wire nc28066;
wire nc28067;
wire nc28068;
wire nc28069;
wire nc28070;
wire nc28071;
wire nc28072;
wire nc28073;
wire nc28074;
wire nc28075;
wire nc28076;
wire nc28077;
wire nc28078;
wire nc28079;
wire nc28080;
wire nc28081;
wire nc28082;
wire nc28083;
wire nc28084;
wire nc28085;
wire nc28086;
wire nc28087;
wire nc28088;
wire nc28089;
wire nc28090;
wire nc28091;
wire nc28092;
wire nc28093;
wire nc28094;
wire nc28095;
wire nc28096;
wire nc28097;
wire nc28098;
wire nc28099;
wire nc28100;
wire nc28101;
wire nc28102;
wire nc28103;
wire nc28104;
wire nc28105;
wire nc28106;
wire nc28107;
wire nc28108;
wire nc28109;
wire nc28110;
wire nc28111;
wire nc28112;
wire nc28113;
wire nc28114;
wire nc28115;
wire nc28116;
wire nc28117;
wire nc28118;
wire nc28119;
wire nc28120;
wire nc28121;
wire nc28122;
wire nc28123;
wire nc28124;
wire nc28125;
wire nc28126;
wire nc28127;
wire nc28128;
wire nc28129;
wire nc28130;
wire nc28131;
wire nc28132;
wire nc28133;
wire nc28134;
wire nc28135;
wire nc28136;
wire nc28137;
wire nc28138;
wire nc28139;
wire nc28140;
wire nc28141;
wire nc28142;
wire nc28143;
wire nc28144;
wire nc28145;
wire nc28146;
wire nc28147;
wire nc28148;
wire nc28149;
wire nc28150;
wire nc28151;
wire nc28152;
wire nc28153;
wire nc28154;
wire nc28155;
wire nc28156;
wire nc28157;
wire nc28158;
wire nc28159;
wire nc28160;
wire nc28161;
wire nc28162;
wire nc28163;
wire nc28164;
wire nc28165;
wire nc28166;
wire nc28167;
wire nc28168;
wire nc28169;
wire nc28170;
wire nc28171;
wire nc28172;
wire nc28173;
wire nc28174;
wire nc28175;
wire nc28176;
wire nc28177;
wire nc28178;
wire nc28179;
wire nc28180;
wire nc28181;
wire nc28182;
wire nc28183;
wire nc28184;
wire nc28185;
wire nc28186;
wire nc28187;
wire nc28188;
wire nc28189;
wire nc28190;
wire nc28191;
wire nc28192;
wire nc28193;
wire nc28194;
wire nc28195;
wire nc28196;
wire nc28197;
wire nc28198;
wire nc28199;
wire nc28200;
wire nc28201;
wire nc28202;
wire nc28203;
wire nc28204;
wire nc28205;
wire nc28206;
wire nc28207;
wire nc28208;
wire nc28209;
wire nc28210;
wire nc28211;
wire nc28212;
wire nc28213;
wire nc28214;
wire nc28215;
wire nc28216;
wire nc28217;
wire nc28218;
wire nc28219;
wire nc28220;
wire nc28221;
wire nc28222;
wire nc28223;
wire nc28224;
wire nc28225;
wire nc28226;
wire nc28227;
wire nc28228;
wire nc28229;
wire nc28230;
wire nc28231;
wire nc28232;
wire nc28233;
wire nc28234;
wire nc28235;
wire nc28236;
wire nc28237;
wire nc28238;
wire nc28239;
wire nc28240;
wire nc28241;
wire nc28242;
wire nc28243;
wire nc28244;
wire nc28245;
wire nc28246;
wire nc28247;
wire nc28248;
wire nc28249;
wire nc28250;
wire nc28251;
wire nc28252;
wire nc28253;
wire nc28254;
wire nc28255;
wire nc28256;
wire nc28257;
wire nc28258;
wire nc28259;
wire nc28260;
wire nc28261;
wire nc28262;
wire nc28263;
wire nc28264;
wire nc28265;
wire nc28266;
wire nc28267;
wire nc28268;
wire nc28269;
wire nc28270;
wire nc28271;
wire nc28272;
wire nc28273;
wire nc28274;
wire nc28275;
wire nc28276;
wire nc28277;
wire nc28278;
wire nc28279;
wire nc28280;
wire nc28281;
wire nc28282;
wire nc28283;
wire nc28284;
wire nc28285;
wire nc28286;
wire nc28287;
wire nc28288;
wire nc28289;
wire nc28290;
wire nc28291;
wire nc28292;
wire nc28293;
wire nc28294;
wire nc28295;
wire nc28296;
wire nc28297;
wire nc28298;
wire nc28299;
wire nc28300;
wire nc28301;
wire nc28302;
wire nc28303;
wire nc28304;
wire nc28305;
wire nc28306;
wire nc28307;
wire nc28308;
wire nc28309;
wire nc28310;
wire nc28311;
wire nc28312;
wire nc28313;
wire nc28314;
wire nc28315;
wire nc28316;
wire nc28317;
wire nc28318;
wire nc28319;
wire nc28320;
wire nc28321;
wire nc28322;
wire nc28323;
wire nc28324;
wire nc28325;
wire nc28326;
wire nc28327;
wire nc28328;
wire nc28329;
wire nc28330;
wire nc28331;
wire nc28332;
wire nc28333;
wire nc28334;
wire nc28335;
wire nc28336;
wire nc28337;
wire nc28338;
wire nc28339;
wire nc28340;
wire nc28341;
wire nc28342;
wire nc28343;
wire nc28344;
wire nc28345;
wire nc28346;
wire nc28347;
wire nc28348;
wire nc28349;
wire nc28350;
wire nc28351;
wire nc28352;
wire nc28353;
wire nc28354;
wire nc28355;
wire nc28356;
wire nc28357;
wire nc28358;
wire nc28359;
wire nc28360;
wire nc28361;
wire nc28362;
wire nc28363;
wire nc28364;
wire nc28365;
wire nc28366;
wire nc28367;
wire nc28368;
wire nc28369;
wire nc28370;
wire nc28371;
wire nc28372;
wire nc28373;
wire nc28374;
wire nc28375;
wire nc28376;
wire nc28377;
wire nc28378;
wire nc28379;
wire nc28380;
wire nc28381;
wire nc28382;
wire nc28383;
wire nc28384;
wire nc28385;
wire nc28386;
wire nc28387;
wire nc28388;
wire nc28389;
wire nc28390;
wire nc28391;
wire nc28392;
wire nc28393;
wire nc28394;
wire nc28395;
wire nc28396;
wire nc28397;
wire nc28398;
wire nc28399;
wire nc28400;
wire nc28401;
wire nc28402;
wire nc28403;
wire nc28404;
wire nc28405;
wire nc28406;
wire nc28407;
wire nc28408;
wire nc28409;
wire nc28410;
wire nc28411;
wire nc28412;
wire nc28413;
wire nc28414;
wire nc28415;
wire nc28416;
wire nc28417;
wire nc28418;
wire nc28419;
wire nc28420;
wire nc28421;
wire nc28422;
wire nc28423;
wire nc28424;
wire nc28425;
wire nc28426;
wire nc28427;
wire nc28428;
wire nc28429;
wire nc28430;
wire nc28431;
wire nc28432;
wire nc28433;
wire nc28434;
wire nc28435;
wire nc28436;
wire nc28437;
wire nc28438;
wire nc28439;
wire nc28440;
wire nc28441;
wire nc28442;
wire nc28443;
wire nc28444;
wire nc28445;
wire nc28446;
wire nc28447;
wire nc28448;
wire nc28449;
wire nc28450;
wire nc28451;
wire nc28452;
wire nc28453;
wire nc28454;
wire nc28455;
wire nc28456;
wire nc28457;
wire nc28458;
wire nc28459;
wire nc28460;
wire nc28461;
wire nc28462;
wire nc28463;
wire nc28464;
wire nc28465;
wire nc28466;
wire nc28467;
wire nc28468;
wire nc28469;
wire nc28470;
wire nc28471;
wire nc28472;
wire nc28473;
wire nc28474;
wire nc28475;
wire nc28476;
wire nc28477;
wire nc28478;
wire nc28479;
wire nc28480;
wire nc28481;
wire nc28482;
wire nc28483;
wire nc28484;
wire nc28485;
wire nc28486;
wire nc28487;
wire nc28488;
wire nc28489;
wire nc28490;
wire nc28491;
wire nc28492;
wire nc28493;
wire nc28494;
wire nc28495;
wire nc28496;
wire nc28497;
wire nc28498;
wire nc28499;
wire nc28500;
wire nc28501;
wire nc28502;
wire nc28503;
wire nc28504;
wire nc28505;
wire nc28506;
wire nc28507;
wire nc28508;
wire nc28509;
wire nc28510;
wire nc28511;
wire nc28512;
wire nc28513;
wire nc28514;
wire nc28515;
wire nc28516;
wire nc28517;
wire nc28518;
wire nc28519;
wire nc28520;
wire nc28521;
wire nc28522;
wire nc28523;
wire nc28524;
wire nc28525;
wire nc28526;
wire nc28527;
wire nc28528;
wire nc28529;
wire nc28530;
wire nc28531;
wire nc28532;
wire nc28533;
wire nc28534;
wire nc28535;
wire nc28536;
wire nc28537;
wire nc28538;
wire nc28539;
wire nc28540;
wire nc28541;
wire nc28542;
wire nc28543;
wire nc28544;
wire nc28545;
wire nc28546;
wire nc28547;
wire nc28548;
wire nc28549;
wire nc28550;
wire nc28551;
wire nc28552;
wire nc28553;
wire nc28554;
wire nc28555;
wire nc28556;
wire nc28557;
wire nc28558;
wire nc28559;
wire nc28560;
wire nc28561;
wire nc28562;
wire nc28563;
wire nc28564;
wire nc28565;
wire nc28566;
wire nc28567;
wire nc28568;
wire nc28569;
wire nc28570;
wire nc28571;
wire nc28572;
wire nc28573;
wire nc28574;
wire nc28575;
wire nc28576;
wire nc28577;
wire nc28578;
wire nc28579;
wire nc28580;
wire nc28581;
wire nc28582;
wire nc28583;
wire nc28584;
wire nc28585;
wire nc28586;
wire nc28587;
wire nc28588;
wire nc28589;
wire nc28590;
wire nc28591;
wire nc28592;
wire nc28593;
wire nc28594;
wire nc28595;
wire nc28596;
wire nc28597;
wire nc28598;
wire nc28599;
wire nc28600;
wire nc28601;
wire nc28602;
wire nc28603;
wire nc28604;
wire nc28605;
wire nc28606;
wire nc28607;
wire nc28608;
wire nc28609;
wire nc28610;
wire nc28611;
wire nc28612;
wire nc28613;
wire nc28614;
wire nc28615;
wire nc28616;
wire nc28617;
wire nc28618;
wire nc28619;
wire nc28620;
wire nc28621;
wire nc28622;
wire nc28623;
wire nc28624;
wire nc28625;
wire nc28626;
wire nc28627;
wire nc28628;
wire nc28629;
wire nc28630;
wire nc28631;
wire nc28632;
wire nc28633;
wire nc28634;
wire nc28635;
wire nc28636;
wire nc28637;
wire nc28638;
wire nc28639;
wire nc28640;
wire nc28641;
wire nc28642;
wire nc28643;
wire nc28644;
wire nc28645;
wire nc28646;
wire nc28647;
wire nc28648;
wire nc28649;
wire nc28650;
wire nc28651;
wire nc28652;
wire nc28653;
wire nc28654;
wire nc28655;
wire nc28656;
wire nc28657;
wire nc28658;
wire nc28659;
wire nc28660;
wire nc28661;
wire nc28662;
wire nc28663;
wire nc28664;
wire nc28665;
wire nc28666;
wire nc28667;
wire nc28668;
wire nc28669;
wire nc28670;
wire nc28671;
wire nc28672;
wire nc28673;
wire nc28674;
wire nc28675;
wire nc28676;
wire nc28677;
wire nc28678;
wire nc28679;
wire nc28680;
wire nc28681;
wire nc28682;
wire nc28683;
wire nc28684;
wire nc28685;
wire nc28686;
wire nc28687;
wire nc28688;
wire nc28689;
wire nc28690;
wire nc28691;
wire nc28692;
wire nc28693;
wire nc28694;
wire nc28695;
wire nc28696;
wire nc28697;
wire nc28698;
wire nc28699;
wire nc28700;
wire nc28701;
wire nc28702;
wire nc28703;
wire nc28704;
wire nc28705;
wire nc28706;
wire nc28707;
wire nc28708;
wire nc28709;
wire nc28710;
wire nc28711;
wire nc28712;
wire nc28713;
wire nc28714;
wire nc28715;
wire nc28716;
wire nc28717;
wire nc28718;
wire nc28719;
wire nc28720;
wire nc28721;
wire nc28722;
wire nc28723;
wire nc28724;
wire nc28725;
wire nc28726;
wire nc28727;
wire nc28728;
wire nc28729;
wire nc28730;
wire nc28731;
wire nc28732;
wire nc28733;
wire nc28734;
wire nc28735;
wire nc28736;
wire nc28737;
wire nc28738;
wire nc28739;
wire nc28740;
wire nc28741;
wire nc28742;
wire nc28743;
wire nc28744;
wire nc28745;
wire nc28746;
wire nc28747;
wire nc28748;
wire nc28749;
wire nc28750;
wire nc28751;
wire nc28752;
wire nc28753;
wire nc28754;
wire nc28755;
wire nc28756;
wire nc28757;
wire nc28758;
wire nc28759;
wire nc28760;
wire nc28761;
wire nc28762;
wire nc28763;
wire nc28764;
wire nc28765;
wire nc28766;
wire nc28767;
wire nc28768;
wire nc28769;
wire nc28770;
wire nc28771;
wire nc28772;
wire nc28773;
wire nc28774;
wire nc28775;
wire nc28776;
wire nc28777;
wire nc28778;
wire nc28779;
wire nc28780;
wire nc28781;
wire nc28782;
wire nc28783;
wire nc28784;
wire nc28785;
wire nc28786;
wire nc28787;
wire nc28788;
wire nc28789;
wire nc28790;
wire nc28791;
wire nc28792;
wire nc28793;
wire nc28794;
wire nc28795;
wire nc28796;
wire nc28797;
wire nc28798;
wire nc28799;
wire nc28800;
wire nc28801;
wire nc28802;
wire nc28803;
wire nc28804;
wire nc28805;
wire nc28806;
wire nc28807;
wire nc28808;
wire nc28809;
wire nc28810;
wire nc28811;
wire nc28812;
wire nc28813;
wire nc28814;
wire nc28815;
wire nc28816;
wire nc28817;
wire nc28818;
wire nc28819;
wire nc28820;
wire nc28821;
wire nc28822;
wire nc28823;
wire nc28824;
wire nc28825;
wire nc28826;
wire nc28827;
wire nc28828;
wire nc28829;
wire nc28830;
wire nc28831;
wire nc28832;
wire nc28833;
wire nc28834;
wire nc28835;
wire nc28836;
wire nc28837;
wire nc28838;
wire nc28839;
wire nc28840;
wire nc28841;
wire nc28842;
wire nc28843;
wire nc28844;
wire nc28845;
wire nc28846;
wire nc28847;
wire nc28848;
wire nc28849;
wire nc28850;
wire nc28851;
wire nc28852;
wire nc28853;
wire nc28854;
wire nc28855;
wire nc28856;
wire nc28857;
wire nc28858;
wire nc28859;
wire nc28860;
wire nc28861;
wire nc28862;
wire nc28863;
wire nc28864;
wire nc28865;
wire nc28866;
wire nc28867;
wire nc28868;
wire nc28869;
wire nc28870;
wire nc28871;
wire nc28872;
wire nc28873;
wire nc28874;
wire nc28875;
wire nc28876;
wire nc28877;
wire nc28878;
wire nc28879;
wire nc28880;
wire nc28881;
wire nc28882;
wire nc28883;
wire nc28884;
wire nc28885;
wire nc28886;
wire nc28887;
wire nc28888;
wire nc28889;
wire nc28890;
wire nc28891;
wire nc28892;
wire nc28893;
wire nc28894;
wire nc28895;
wire nc28896;
wire nc28897;
wire nc28898;
wire nc28899;
wire nc28900;
wire nc28901;
wire nc28902;
wire nc28903;
wire nc28904;
wire nc28905;
wire nc28906;
wire nc28907;
wire nc28908;
wire nc28909;
wire nc28910;
wire nc28911;
wire nc28912;
wire nc28913;
wire nc28914;
wire nc28915;
wire nc28916;
wire nc28917;
wire nc28918;
wire nc28919;
wire nc28920;
wire nc28921;
wire nc28922;
wire nc28923;
wire nc28924;
wire nc28925;
wire nc28926;
wire nc28927;
wire nc28928;
wire nc28929;
wire nc28930;
wire nc28931;
wire nc28932;
wire nc28933;
wire nc28934;
wire nc28935;
wire nc28936;
wire nc28937;
wire nc28938;
wire nc28939;
wire nc28940;
wire nc28941;
wire nc28942;
wire nc28943;
wire nc28944;
wire nc28945;
wire nc28946;
wire nc28947;
wire nc28948;
wire nc28949;
wire nc28950;
wire nc28951;
wire nc28952;
wire nc28953;
wire nc28954;
wire nc28955;
wire nc28956;
wire nc28957;
wire nc28958;
wire nc28959;
wire nc28960;
wire nc28961;
wire nc28962;
wire nc28963;
wire nc28964;
wire nc28965;
wire nc28966;
wire nc28967;
wire nc28968;
wire nc28969;
wire nc28970;
wire nc28971;
wire nc28972;
wire nc28973;
wire nc28974;
wire nc28975;
wire nc28976;
wire nc28977;
wire nc28978;
wire nc28979;
wire nc28980;
wire nc28981;
wire nc28982;
wire nc28983;
wire nc28984;
wire nc28985;
wire nc28986;
wire nc28987;
wire nc28988;
wire nc28989;
wire nc28990;
wire nc28991;
wire nc28992;
wire nc28993;
wire nc28994;
wire nc28995;
wire nc28996;
wire nc28997;
wire nc28998;
wire nc28999;
wire nc29000;
wire nc29001;
wire nc29002;
wire nc29003;
wire nc29004;
wire nc29005;
wire nc29006;
wire nc29007;
wire nc29008;
wire nc29009;
wire nc29010;
wire nc29011;
wire nc29012;
wire nc29013;
wire nc29014;
wire nc29015;
wire nc29016;
wire nc29017;
wire nc29018;
wire nc29019;
wire nc29020;
wire nc29021;
wire nc29022;
wire nc29023;
wire nc29024;
wire nc29025;
wire nc29026;
wire nc29027;
wire nc29028;
wire nc29029;
wire nc29030;
wire nc29031;
wire nc29032;
wire nc29033;
wire nc29034;
wire nc29035;
wire nc29036;
wire nc29037;
wire nc29038;
wire nc29039;
wire nc29040;
wire nc29041;
wire nc29042;
wire nc29043;
wire nc29044;
wire nc29045;
wire nc29046;
wire nc29047;
wire nc29048;
wire nc29049;
wire nc29050;
wire nc29051;
wire nc29052;
wire nc29053;
wire nc29054;
wire nc29055;
wire nc29056;
wire nc29057;
wire nc29058;
wire nc29059;
wire nc29060;
wire nc29061;
wire nc29062;
wire nc29063;
wire nc29064;
wire nc29065;
wire nc29066;
wire nc29067;
wire nc29068;
wire nc29069;
wire nc29070;
wire nc29071;
wire nc29072;
wire nc29073;
wire nc29074;
wire nc29075;
wire nc29076;
wire nc29077;
wire nc29078;
wire nc29079;
wire nc29080;
wire nc29081;
wire nc29082;
wire nc29083;
wire nc29084;
wire nc29085;
wire nc29086;
wire nc29087;
wire nc29088;
wire nc29089;
wire nc29090;
wire nc29091;
wire nc29092;
wire nc29093;
wire nc29094;
wire nc29095;
wire nc29096;
wire nc29097;
wire nc29098;
wire nc29099;
wire nc29100;
wire nc29101;
wire nc29102;
wire nc29103;
wire nc29104;
wire nc29105;
wire nc29106;
wire nc29107;
wire nc29108;
wire nc29109;
wire nc29110;
wire nc29111;
wire nc29112;
wire nc29113;
wire nc29114;
wire nc29115;
wire nc29116;
wire nc29117;
wire nc29118;
wire nc29119;
wire nc29120;
wire nc29121;
wire nc29122;
wire nc29123;
wire nc29124;
wire nc29125;
wire nc29126;
wire nc29127;
wire nc29128;
wire nc29129;
wire nc29130;
wire nc29131;
wire nc29132;
wire nc29133;
wire nc29134;
wire nc29135;
wire nc29136;
wire nc29137;
wire nc29138;
wire nc29139;
wire nc29140;
wire nc29141;
wire nc29142;
wire nc29143;
wire nc29144;
wire nc29145;
wire nc29146;
wire nc29147;
wire nc29148;
wire nc29149;
wire nc29150;
wire nc29151;
wire nc29152;
wire nc29153;
wire nc29154;
wire nc29155;
wire nc29156;
wire nc29157;
wire nc29158;
wire nc29159;
wire nc29160;
wire nc29161;
wire nc29162;
wire nc29163;
wire nc29164;
wire nc29165;
wire nc29166;
wire nc29167;
wire nc29168;
wire nc29169;
wire nc29170;
wire nc29171;
wire nc29172;
wire nc29173;
wire nc29174;
wire nc29175;
wire nc29176;
wire nc29177;
wire nc29178;
wire nc29179;
wire nc29180;
wire nc29181;
wire nc29182;
wire nc29183;
wire nc29184;
wire nc29185;
wire nc29186;
wire nc29187;
wire nc29188;
wire nc29189;
wire nc29190;
wire nc29191;
wire nc29192;
wire nc29193;
wire nc29194;
wire nc29195;
wire nc29196;
wire nc29197;
wire nc29198;
wire nc29199;
wire nc29200;
wire nc29201;
wire nc29202;
wire nc29203;
wire nc29204;
wire nc29205;
wire nc29206;
wire nc29207;
wire nc29208;
wire nc29209;
wire nc29210;
wire nc29211;
wire nc29212;
wire nc29213;
wire nc29214;
wire nc29215;
wire nc29216;
wire nc29217;
wire nc29218;
wire nc29219;
wire nc29220;
wire nc29221;
wire nc29222;
wire nc29223;
wire nc29224;
wire nc29225;
wire nc29226;
wire nc29227;
wire nc29228;
wire nc29229;
wire nc29230;
wire nc29231;
wire nc29232;
wire nc29233;
wire nc29234;
wire nc29235;
wire nc29236;
wire nc29237;
wire nc29238;
wire nc29239;
wire nc29240;
wire nc29241;
wire nc29242;
wire nc29243;
wire nc29244;
wire nc29245;
wire nc29246;
wire nc29247;
wire nc29248;
wire nc29249;
wire nc29250;
wire nc29251;
wire nc29252;
wire nc29253;
wire nc29254;
wire nc29255;
wire nc29256;
wire nc29257;
wire nc29258;
wire nc29259;
wire nc29260;
wire nc29261;
wire nc29262;
wire nc29263;
wire nc29264;
wire nc29265;
wire nc29266;
wire nc29267;
wire nc29268;
wire nc29269;
wire nc29270;
wire nc29271;
wire nc29272;
wire nc29273;
wire nc29274;
wire nc29275;
wire nc29276;
wire nc29277;
wire nc29278;
wire nc29279;
wire nc29280;
wire nc29281;
wire nc29282;
wire nc29283;
wire nc29284;
wire nc29285;
wire nc29286;
wire nc29287;
wire nc29288;
wire nc29289;
wire nc29290;
wire nc29291;
wire nc29292;
wire nc29293;
wire nc29294;
wire nc29295;
wire nc29296;
wire nc29297;
wire nc29298;
wire nc29299;
wire nc29300;
wire nc29301;
wire nc29302;
wire nc29303;
wire nc29304;
wire nc29305;
wire nc29306;
wire nc29307;
wire nc29308;
wire nc29309;
wire nc29310;
wire nc29311;
wire nc29312;
wire nc29313;
wire nc29314;
wire nc29315;
wire nc29316;
wire nc29317;
wire nc29318;
wire nc29319;
wire nc29320;
wire nc29321;
wire nc29322;
wire nc29323;
wire nc29324;
wire nc29325;
wire nc29326;
wire nc29327;
wire nc29328;
wire nc29329;
wire nc29330;
wire nc29331;
wire nc29332;
wire nc29333;
wire nc29334;
wire nc29335;
wire nc29336;
wire nc29337;
wire nc29338;
wire nc29339;
wire nc29340;
wire nc29341;
wire nc29342;
wire nc29343;
wire nc29344;
wire nc29345;
wire nc29346;
wire nc29347;
wire nc29348;
wire nc29349;
wire nc29350;
wire nc29351;
wire nc29352;
wire nc29353;
wire nc29354;
wire nc29355;
wire nc29356;
wire nc29357;
wire nc29358;
wire nc29359;
wire nc29360;
wire nc29361;
wire nc29362;
wire nc29363;
wire nc29364;
wire nc29365;
wire nc29366;
wire nc29367;
wire nc29368;
wire nc29369;
wire nc29370;
wire nc29371;
wire nc29372;
wire nc29373;
wire nc29374;
wire nc29375;
wire nc29376;
wire nc29377;
wire nc29378;
wire nc29379;
wire nc29380;
wire nc29381;
wire nc29382;
wire nc29383;
wire nc29384;
wire nc29385;
wire nc29386;
wire nc29387;
wire nc29388;
wire nc29389;
wire nc29390;
wire nc29391;
wire nc29392;
wire nc29393;
wire nc29394;
wire nc29395;
wire nc29396;
wire nc29397;
wire nc29398;
wire nc29399;
wire nc29400;
wire nc29401;
wire nc29402;
wire nc29403;
wire nc29404;
wire nc29405;
wire nc29406;
wire nc29407;
wire nc29408;
wire nc29409;
wire nc29410;
wire nc29411;
wire nc29412;
wire nc29413;
wire nc29414;
wire nc29415;
wire nc29416;
wire nc29417;
wire nc29418;
wire nc29419;
wire nc29420;
wire nc29421;
wire nc29422;
wire nc29423;
wire nc29424;
wire nc29425;
wire nc29426;
wire nc29427;
wire nc29428;
wire nc29429;
wire nc29430;
wire nc29431;
wire nc29432;
wire nc29433;
wire nc29434;
wire nc29435;
wire nc29436;
wire nc29437;
wire nc29438;
wire nc29439;
wire nc29440;
wire nc29441;
wire nc29442;
wire nc29443;
wire nc29444;
wire nc29445;
wire nc29446;
wire nc29447;
wire nc29448;
wire nc29449;
wire nc29450;
wire nc29451;
wire nc29452;
wire nc29453;
wire nc29454;
wire nc29455;
wire nc29456;
wire nc29457;
wire nc29458;
wire nc29459;
wire nc29460;
wire nc29461;
wire nc29462;
wire nc29463;
wire nc29464;
wire nc29465;
wire nc29466;
wire nc29467;
wire nc29468;
wire nc29469;
wire nc29470;
wire nc29471;
wire nc29472;
wire nc29473;
wire nc29474;
wire nc29475;
wire nc29476;
wire nc29477;
wire nc29478;
wire nc29479;
wire nc29480;
wire nc29481;
wire nc29482;
wire nc29483;
wire nc29484;
wire nc29485;
wire nc29486;
wire nc29487;
wire nc29488;
wire nc29489;
wire nc29490;
wire nc29491;
wire nc29492;
wire nc29493;
wire nc29494;
wire nc29495;
wire nc29496;
wire nc29497;
wire nc29498;
wire nc29499;
wire nc29500;
wire nc29501;
wire nc29502;
wire nc29503;
wire nc29504;
wire nc29505;
wire nc29506;
wire nc29507;
wire nc29508;
wire nc29509;
wire nc29510;
wire nc29511;
wire nc29512;
wire nc29513;
wire nc29514;
wire nc29515;
wire nc29516;
wire nc29517;
wire nc29518;
wire nc29519;
wire nc29520;
wire nc29521;
wire nc29522;
wire nc29523;
wire nc29524;
wire nc29525;
wire nc29526;
wire nc29527;
wire nc29528;
wire nc29529;
wire nc29530;
wire nc29531;
wire nc29532;
wire nc29533;
wire nc29534;
wire nc29535;
wire nc29536;
wire nc29537;
wire nc29538;
wire nc29539;
wire nc29540;
wire nc29541;
wire nc29542;
wire nc29543;
wire nc29544;
wire nc29545;
wire nc29546;
wire nc29547;
wire nc29548;
wire nc29549;
wire nc29550;
wire nc29551;
wire nc29552;
wire nc29553;
wire nc29554;
wire nc29555;
wire nc29556;
wire nc29557;
wire nc29558;
wire nc29559;
wire nc29560;
wire nc29561;
wire nc29562;
wire nc29563;
wire nc29564;
wire nc29565;
wire nc29566;
wire nc29567;
wire nc29568;
wire nc29569;
wire nc29570;
wire nc29571;
wire nc29572;
wire nc29573;
wire nc29574;
wire nc29575;
wire nc29576;
wire nc29577;
wire nc29578;
wire nc29579;
wire nc29580;
wire nc29581;
wire nc29582;
wire nc29583;
wire nc29584;
wire nc29585;
wire nc29586;
wire nc29587;
wire nc29588;
wire nc29589;
wire nc29590;
wire nc29591;
wire nc29592;
wire nc29593;
wire nc29594;
wire nc29595;
wire nc29596;
wire nc29597;
wire nc29598;
wire nc29599;
wire nc29600;
wire nc29601;
wire nc29602;
wire nc29603;
wire nc29604;
wire nc29605;
wire nc29606;
wire nc29607;
wire nc29608;
wire nc29609;
wire nc29610;
wire nc29611;
wire nc29612;
wire nc29613;
wire nc29614;
wire nc29615;
wire nc29616;
wire nc29617;
wire nc29618;
wire nc29619;
wire nc29620;
wire nc29621;
wire nc29622;
wire nc29623;
wire nc29624;
wire nc29625;
wire nc29626;
wire nc29627;
wire nc29628;
wire nc29629;
wire nc29630;
wire nc29631;
wire nc29632;
wire nc29633;
wire nc29634;
wire nc29635;
wire nc29636;
wire nc29637;
wire nc29638;
wire nc29639;
wire nc29640;
wire nc29641;
wire nc29642;
wire nc29643;
wire nc29644;
wire nc29645;
wire nc29646;
wire nc29647;
wire nc29648;
wire nc29649;
wire nc29650;
wire nc29651;
wire nc29652;
wire nc29653;
wire nc29654;
wire nc29655;
wire nc29656;
wire nc29657;
wire nc29658;
wire nc29659;
wire nc29660;
wire nc29661;
wire nc29662;
wire nc29663;
wire nc29664;
wire nc29665;
wire nc29666;
wire nc29667;
wire nc29668;
wire nc29669;
wire nc29670;
wire nc29671;
wire nc29672;
wire nc29673;
wire nc29674;
wire nc29675;
wire nc29676;
wire nc29677;
wire nc29678;
wire nc29679;
wire nc29680;
wire nc29681;
wire nc29682;
wire nc29683;
wire nc29684;
wire nc29685;
wire nc29686;
wire nc29687;
wire nc29688;
wire nc29689;
wire nc29690;
wire nc29691;
wire nc29692;
wire nc29693;
wire nc29694;
wire nc29695;
wire nc29696;
wire nc29697;
wire nc29698;
wire nc29699;
wire nc29700;
wire nc29701;
wire nc29702;
wire nc29703;
wire nc29704;
wire nc29705;
wire nc29706;
wire nc29707;
wire nc29708;
wire nc29709;
wire nc29710;
wire nc29711;
wire nc29712;
wire nc29713;
wire nc29714;
wire nc29715;
wire nc29716;
wire nc29717;
wire nc29718;
wire nc29719;
wire nc29720;
wire nc29721;
wire nc29722;
wire nc29723;
wire nc29724;
wire nc29725;
wire nc29726;
wire nc29727;
wire nc29728;
wire nc29729;
wire nc29730;
wire nc29731;
wire nc29732;
wire nc29733;
wire nc29734;
wire nc29735;
wire nc29736;
wire nc29737;
wire nc29738;
wire nc29739;
wire nc29740;
wire nc29741;
wire nc29742;
wire nc29743;
wire nc29744;
wire nc29745;
wire nc29746;
wire nc29747;
wire nc29748;
wire nc29749;
wire nc29750;
wire nc29751;
wire nc29752;
wire nc29753;
wire nc29754;
wire nc29755;
wire nc29756;
wire nc29757;
wire nc29758;
wire nc29759;
wire nc29760;
wire nc29761;
wire nc29762;
wire nc29763;
wire nc29764;
wire nc29765;
wire nc29766;
wire nc29767;
wire nc29768;
wire nc29769;
wire nc29770;
wire nc29771;
wire nc29772;
wire nc29773;
wire nc29774;
wire nc29775;
wire nc29776;
wire nc29777;
wire nc29778;
wire nc29779;
wire nc29780;
wire nc29781;
wire nc29782;
wire nc29783;
wire nc29784;
wire nc29785;
wire nc29786;
wire nc29787;
wire nc29788;
wire nc29789;
wire nc29790;
wire nc29791;
wire nc29792;
wire nc29793;
wire nc29794;
wire nc29795;
wire nc29796;
wire nc29797;
wire nc29798;
wire nc29799;
wire nc29800;
wire nc29801;
wire nc29802;
wire nc29803;
wire nc29804;
wire nc29805;
wire nc29806;
wire nc29807;
wire nc29808;
wire nc29809;
wire nc29810;
wire nc29811;
wire nc29812;
wire nc29813;
wire nc29814;
wire nc29815;
wire nc29816;
wire nc29817;
wire nc29818;
wire nc29819;
wire nc29820;
wire nc29821;
wire nc29822;
wire nc29823;
wire nc29824;
wire nc29825;
wire nc29826;
wire nc29827;
wire nc29828;
wire nc29829;
wire nc29830;
wire nc29831;
wire nc29832;
wire nc29833;
wire nc29834;
wire nc29835;
wire nc29836;
wire nc29837;
wire nc29838;
wire nc29839;
wire nc29840;
wire nc29841;
wire nc29842;
wire nc29843;
wire nc29844;
wire nc29845;
wire nc29846;
wire nc29847;
wire nc29848;
wire nc29849;
wire nc29850;
wire nc29851;
wire nc29852;
wire nc29853;
wire nc29854;
wire nc29855;
wire nc29856;
wire nc29857;
wire nc29858;
wire nc29859;
wire nc29860;
wire nc29861;
wire nc29862;
wire nc29863;
wire nc29864;
wire nc29865;
wire nc29866;
wire nc29867;
wire nc29868;
wire nc29869;
wire nc29870;
wire nc29871;
wire nc29872;
wire nc29873;
wire nc29874;
wire nc29875;
wire nc29876;
wire nc29877;
wire nc29878;
wire nc29879;
wire nc29880;
wire nc29881;
wire nc29882;
wire nc29883;
wire nc29884;
wire nc29885;
wire nc29886;
wire nc29887;
wire nc29888;
wire nc29889;
wire nc29890;
wire nc29891;
wire nc29892;
wire nc29893;
wire nc29894;
wire nc29895;
wire nc29896;
wire nc29897;
wire nc29898;
wire nc29899;
wire nc29900;
wire nc29901;
wire nc29902;
wire nc29903;
wire nc29904;
wire nc29905;
wire nc29906;
wire nc29907;
wire nc29908;
wire nc29909;
wire nc29910;
wire nc29911;
wire nc29912;
wire nc29913;
wire nc29914;
wire nc29915;
wire nc29916;
wire nc29917;
wire nc29918;
wire nc29919;
wire nc29920;
wire nc29921;
wire nc29922;
wire nc29923;
wire nc29924;
wire nc29925;
wire nc29926;
wire nc29927;
wire nc29928;
wire nc29929;
wire nc29930;
wire nc29931;
wire nc29932;
wire nc29933;
wire nc29934;
wire nc29935;
wire nc29936;
wire nc29937;
wire nc29938;
wire nc29939;
wire nc29940;
wire nc29941;
wire nc29942;
wire nc29943;
wire nc29944;
wire nc29945;
wire nc29946;
wire nc29947;
wire nc29948;
wire nc29949;
wire nc29950;
wire nc29951;
wire nc29952;
wire nc29953;
wire nc29954;
wire nc29955;
wire nc29956;
wire nc29957;
wire nc29958;
wire nc29959;
wire nc29960;
wire nc29961;
wire nc29962;
wire nc29963;
wire nc29964;
wire nc29965;
wire nc29966;
wire nc29967;
wire nc29968;
wire nc29969;
wire nc29970;
wire nc29971;
wire nc29972;
wire nc29973;
wire nc29974;
wire nc29975;
wire nc29976;
wire nc29977;
wire nc29978;
wire nc29979;
wire nc29980;
wire nc29981;
wire nc29982;
wire nc29983;
wire nc29984;
wire nc29985;
wire nc29986;
wire nc29987;
wire nc29988;
wire nc29989;
wire nc29990;
wire nc29991;
wire nc29992;
wire nc29993;
wire nc29994;
wire nc29995;
wire nc29996;
wire nc29997;
wire nc29998;
wire nc29999;
wire nc30000;
wire nc30001;
wire nc30002;
wire nc30003;
wire nc30004;
wire nc30005;
wire nc30006;
wire nc30007;
wire nc30008;
wire nc30009;
wire nc30010;
wire nc30011;
wire nc30012;
wire nc30013;
wire nc30014;
wire nc30015;
wire nc30016;
wire nc30017;
wire nc30018;
wire nc30019;
wire nc30020;
wire nc30021;
wire nc30022;
wire nc30023;
wire nc30024;
wire nc30025;
wire nc30026;
wire nc30027;
wire nc30028;
wire nc30029;
wire nc30030;
wire nc30031;
wire nc30032;
wire nc30033;
wire nc30034;
wire nc30035;
wire nc30036;
wire nc30037;
wire nc30038;
wire nc30039;
wire nc30040;
wire nc30041;
wire nc30042;
wire nc30043;
wire nc30044;
wire nc30045;
wire nc30046;
wire nc30047;
wire nc30048;
wire nc30049;
wire nc30050;
wire nc30051;
wire nc30052;
wire nc30053;
wire nc30054;
wire nc30055;
wire nc30056;
wire nc30057;
wire nc30058;
wire nc30059;
wire nc30060;
wire nc30061;
wire nc30062;
wire nc30063;
wire nc30064;
wire nc30065;
wire nc30066;
wire nc30067;
wire nc30068;
wire nc30069;
wire nc30070;
wire nc30071;
wire nc30072;
wire nc30073;
wire nc30074;
wire nc30075;
wire nc30076;
wire nc30077;
wire nc30078;
wire nc30079;
wire nc30080;
wire nc30081;
wire nc30082;
wire nc30083;
wire nc30084;
wire nc30085;
wire nc30086;
wire nc30087;
wire nc30088;
wire nc30089;
wire nc30090;
wire nc30091;
wire nc30092;
wire nc30093;
wire nc30094;
wire nc30095;
wire nc30096;
wire nc30097;
wire nc30098;
wire nc30099;
wire nc30100;
wire nc30101;
wire nc30102;
wire nc30103;
wire nc30104;
wire nc30105;
wire nc30106;
wire nc30107;
wire nc30108;
wire nc30109;
wire nc30110;
wire nc30111;
wire nc30112;
wire nc30113;
wire nc30114;
wire nc30115;
wire nc30116;
wire nc30117;
wire nc30118;
wire nc30119;
wire nc30120;
wire nc30121;
wire nc30122;
wire nc30123;
wire nc30124;
wire nc30125;
wire nc30126;
wire nc30127;
wire nc30128;
wire nc30129;
wire nc30130;
wire nc30131;
wire nc30132;
wire nc30133;
wire nc30134;
wire nc30135;
wire nc30136;
wire nc30137;
wire nc30138;
wire nc30139;
wire nc30140;
wire nc30141;
wire nc30142;
wire nc30143;
wire nc30144;
wire nc30145;
wire nc30146;
wire nc30147;
wire nc30148;
wire nc30149;
wire nc30150;
wire nc30151;
wire nc30152;
wire nc30153;
wire nc30154;
wire nc30155;
wire nc30156;
wire nc30157;
wire nc30158;
wire nc30159;
wire nc30160;
wire nc30161;
wire nc30162;
wire nc30163;
wire nc30164;
wire nc30165;
wire nc30166;
wire nc30167;
wire nc30168;
wire nc30169;
wire nc30170;
wire nc30171;
wire nc30172;
wire nc30173;
wire nc30174;
wire nc30175;
wire nc30176;
wire nc30177;
wire nc30178;
wire nc30179;
wire nc30180;
wire nc30181;
wire nc30182;
wire nc30183;
wire nc30184;
wire nc30185;
wire nc30186;
wire nc30187;
wire nc30188;
wire nc30189;
wire nc30190;
wire nc30191;
wire nc30192;
wire nc30193;
wire nc30194;
wire nc30195;
wire nc30196;
wire nc30197;
wire nc30198;
wire nc30199;
wire nc30200;
wire nc30201;
wire nc30202;
wire nc30203;
wire nc30204;
wire nc30205;
wire nc30206;
wire nc30207;
wire nc30208;
wire nc30209;
wire nc30210;
wire nc30211;
wire nc30212;
wire nc30213;
wire nc30214;
wire nc30215;
wire nc30216;
wire nc30217;
wire nc30218;
wire nc30219;
wire nc30220;
wire nc30221;
wire nc30222;
wire nc30223;
wire nc30224;
wire nc30225;
wire nc30226;
wire nc30227;
wire nc30228;
wire nc30229;
wire nc30230;
wire nc30231;
wire nc30232;
wire nc30233;
wire nc30234;
wire nc30235;
wire nc30236;
wire nc30237;
wire nc30238;
wire nc30239;
wire nc30240;
wire nc30241;
wire nc30242;
wire nc30243;
wire nc30244;
wire nc30245;
wire nc30246;
wire nc30247;
wire nc30248;
wire nc30249;
wire nc30250;
wire nc30251;
wire nc30252;
wire nc30253;
wire nc30254;
wire nc30255;
wire nc30256;
wire nc30257;
wire nc30258;
wire nc30259;
wire nc30260;
wire nc30261;
wire nc30262;
wire nc30263;
wire nc30264;
wire nc30265;
wire nc30266;
wire nc30267;
wire nc30268;
wire nc30269;
wire nc30270;
wire nc30271;
wire nc30272;
wire nc30273;
wire nc30274;
wire nc30275;
wire nc30276;
wire nc30277;
wire nc30278;
wire nc30279;
wire nc30280;
wire nc30281;
wire nc30282;
wire nc30283;
wire nc30284;
wire nc30285;
wire nc30286;
wire nc30287;
wire nc30288;
wire nc30289;
wire nc30290;
wire nc30291;
wire nc30292;
wire nc30293;
wire nc30294;
wire nc30295;
wire nc30296;
wire nc30297;
wire nc30298;
wire nc30299;
wire nc30300;
wire nc30301;
wire nc30302;
wire nc30303;
wire nc30304;
wire nc30305;
wire nc30306;
wire nc30307;
wire nc30308;
wire nc30309;
wire nc30310;
wire nc30311;
wire nc30312;
wire nc30313;
wire nc30314;
wire nc30315;
wire nc30316;
wire nc30317;
wire nc30318;
wire nc30319;
wire nc30320;
wire nc30321;
wire nc30322;
wire nc30323;
wire nc30324;
wire nc30325;
wire nc30326;
wire nc30327;
wire nc30328;
wire nc30329;
wire nc30330;
wire nc30331;
wire nc30332;
wire nc30333;
wire nc30334;
wire nc30335;
wire nc30336;
wire nc30337;
wire nc30338;
wire nc30339;
wire nc30340;
wire nc30341;
wire nc30342;
wire nc30343;
wire nc30344;
wire nc30345;
wire nc30346;
wire nc30347;
wire nc30348;
wire nc30349;
wire nc30350;
wire nc30351;
wire nc30352;
wire nc30353;
wire nc30354;
wire nc30355;
wire nc30356;
wire nc30357;
wire nc30358;
wire nc30359;
wire nc30360;
wire nc30361;
wire nc30362;
wire nc30363;
wire nc30364;
wire nc30365;
wire nc30366;
wire nc30367;
wire nc30368;
wire nc30369;
wire nc30370;
wire nc30371;
wire nc30372;
wire nc30373;
wire nc30374;
wire nc30375;
wire nc30376;
wire nc30377;
wire nc30378;
wire nc30379;
wire nc30380;
wire nc30381;
wire nc30382;
wire nc30383;
wire nc30384;
wire nc30385;
wire nc30386;
wire nc30387;
wire nc30388;
wire nc30389;
wire nc30390;
wire nc30391;
wire nc30392;
wire nc30393;
wire nc30394;
wire nc30395;
wire nc30396;
wire nc30397;
wire nc30398;
wire nc30399;
wire nc30400;
wire nc30401;
wire nc30402;
wire nc30403;
wire nc30404;
wire nc30405;
wire nc30406;
wire nc30407;
wire nc30408;
wire nc30409;
wire nc30410;
wire nc30411;
wire nc30412;
wire nc30413;
wire nc30414;
wire nc30415;
wire nc30416;
wire nc30417;
wire nc30418;
wire nc30419;
wire nc30420;
wire nc30421;
wire nc30422;
wire nc30423;
wire nc30424;
wire nc30425;
wire nc30426;
wire nc30427;
wire nc30428;
wire nc30429;
wire nc30430;
wire nc30431;
wire nc30432;
wire nc30433;
wire nc30434;
wire nc30435;
wire nc30436;
wire nc30437;
wire nc30438;
wire nc30439;
wire nc30440;
wire nc30441;
wire nc30442;
wire nc30443;
wire nc30444;
wire nc30445;
wire nc30446;
wire nc30447;
wire nc30448;
wire nc30449;
wire nc30450;
wire nc30451;
wire nc30452;
wire nc30453;
wire nc30454;
wire nc30455;
wire nc30456;
wire nc30457;
wire nc30458;
wire nc30459;
wire nc30460;
wire nc30461;
wire nc30462;
wire nc30463;
wire nc30464;
wire nc30465;
wire nc30466;
wire nc30467;
wire nc30468;
wire nc30469;
wire nc30470;
wire nc30471;
wire nc30472;
wire nc30473;
wire nc30474;
wire nc30475;
wire nc30476;
wire nc30477;
wire nc30478;
wire nc30479;
wire nc30480;
wire nc30481;
wire nc30482;
wire nc30483;
wire nc30484;
wire nc30485;
wire nc30486;
wire nc30487;
wire nc30488;
wire nc30489;
wire nc30490;
wire nc30491;
wire nc30492;
wire nc30493;
wire nc30494;
wire nc30495;
wire nc30496;
wire nc30497;
wire nc30498;
wire nc30499;
wire nc30500;
wire nc30501;
wire nc30502;
wire nc30503;
wire nc30504;
wire nc30505;
wire nc30506;
wire nc30507;
wire nc30508;
wire nc30509;
wire nc30510;
wire nc30511;
wire nc30512;
wire nc30513;
wire nc30514;
wire nc30515;
wire nc30516;
wire nc30517;
wire nc30518;
wire nc30519;
wire nc30520;
wire nc30521;
wire nc30522;
wire nc30523;
wire nc30524;
wire nc30525;
wire nc30526;
wire nc30527;
wire nc30528;
wire nc30529;
wire nc30530;
wire nc30531;
wire nc30532;
wire nc30533;
wire nc30534;
wire nc30535;
wire nc30536;
wire nc30537;
wire nc30538;
wire nc30539;
wire nc30540;
wire nc30541;
wire nc30542;
wire nc30543;
wire nc30544;
wire nc30545;
wire nc30546;
wire nc30547;
wire nc30548;
wire nc30549;
wire nc30550;
wire nc30551;
wire nc30552;
wire nc30553;
wire nc30554;
wire nc30555;
wire nc30556;
wire nc30557;
wire nc30558;
wire nc30559;
wire nc30560;
wire nc30561;
wire nc30562;
wire nc30563;
wire nc30564;
wire nc30565;
wire nc30566;
wire nc30567;
wire nc30568;
wire nc30569;
wire nc30570;
wire nc30571;
wire nc30572;
wire nc30573;
wire nc30574;
wire nc30575;
wire nc30576;
wire nc30577;
wire nc30578;
wire nc30579;
wire nc30580;
wire nc30581;
wire nc30582;
wire nc30583;
wire nc30584;
wire nc30585;
wire nc30586;
wire nc30587;
wire nc30588;
wire nc30589;
wire nc30590;
wire nc30591;
wire nc30592;
wire nc30593;
wire nc30594;
wire nc30595;
wire nc30596;
wire nc30597;
wire nc30598;
wire nc30599;
wire nc30600;
wire nc30601;
wire nc30602;
wire nc30603;
wire nc30604;
wire nc30605;
wire nc30606;
wire nc30607;
wire nc30608;
wire nc30609;
wire nc30610;
wire nc30611;
wire nc30612;
wire nc30613;
wire nc30614;
wire nc30615;
wire nc30616;
wire nc30617;
wire nc30618;
wire nc30619;
wire nc30620;
wire nc30621;
wire nc30622;
wire nc30623;
wire nc30624;
wire nc30625;
wire nc30626;
wire nc30627;
wire nc30628;
wire nc30629;
wire nc30630;
wire nc30631;
wire nc30632;
wire nc30633;
wire nc30634;
wire nc30635;
wire nc30636;
wire nc30637;
wire nc30638;
wire nc30639;
wire nc30640;
wire nc30641;
wire nc30642;
wire nc30643;
wire nc30644;
wire nc30645;
wire nc30646;
wire nc30647;
wire nc30648;
wire nc30649;
wire nc30650;
wire nc30651;
wire nc30652;
wire nc30653;
wire nc30654;
wire nc30655;
wire nc30656;
wire nc30657;
wire nc30658;
wire nc30659;
wire nc30660;
wire nc30661;
wire nc30662;
wire nc30663;
wire nc30664;
wire nc30665;
wire nc30666;
wire nc30667;
wire nc30668;
wire nc30669;
wire nc30670;
wire nc30671;
wire nc30672;
wire nc30673;
wire nc30674;
wire nc30675;
wire nc30676;
wire nc30677;
wire nc30678;
wire nc30679;
wire nc30680;
wire nc30681;
wire nc30682;
wire nc30683;
wire nc30684;
wire nc30685;
wire nc30686;
wire nc30687;
wire nc30688;
wire nc30689;
wire nc30690;
wire nc30691;
wire nc30692;
wire nc30693;
wire nc30694;
wire nc30695;
wire nc30696;
wire nc30697;
wire nc30698;
wire nc30699;
wire nc30700;
wire nc30701;
wire nc30702;
wire nc30703;
wire nc30704;
wire nc30705;
wire nc30706;
wire nc30707;
wire nc30708;
wire nc30709;
wire nc30710;
wire nc30711;
wire nc30712;
wire nc30713;
wire nc30714;
wire nc30715;
wire nc30716;
wire nc30717;
wire nc30718;
wire nc30719;
wire nc30720;
wire nc30721;
wire nc30722;
wire nc30723;
wire nc30724;
wire nc30725;
wire nc30726;
wire nc30727;
wire nc30728;
wire nc30729;
wire nc30730;
wire nc30731;
wire nc30732;
wire nc30733;
wire nc30734;
wire nc30735;
wire nc30736;
wire nc30737;
wire nc30738;
wire nc30739;
wire nc30740;
wire nc30741;
wire nc30742;
wire nc30743;
wire nc30744;
wire nc30745;
wire nc30746;
wire nc30747;
wire nc30748;
wire nc30749;
wire nc30750;
wire nc30751;
wire nc30752;
wire nc30753;
wire nc30754;
wire nc30755;
wire nc30756;
wire nc30757;
wire nc30758;
wire nc30759;
wire nc30760;
wire nc30761;
wire nc30762;
wire nc30763;
wire nc30764;
wire nc30765;
wire nc30766;
wire nc30767;
wire nc30768;
wire nc30769;
wire nc30770;
wire nc30771;
wire nc30772;
wire nc30773;
wire nc30774;
wire nc30775;
wire nc30776;
wire nc30777;
wire nc30778;
wire nc30779;
wire nc30780;
wire nc30781;
wire nc30782;
wire nc30783;
wire nc30784;
wire nc30785;
wire nc30786;
wire nc30787;
wire nc30788;
wire nc30789;
wire nc30790;
wire nc30791;
wire nc30792;
wire nc30793;
wire nc30794;
wire nc30795;
wire nc30796;
wire nc30797;
wire nc30798;
wire nc30799;
wire nc30800;
wire nc30801;
wire nc30802;
wire nc30803;
wire nc30804;
wire nc30805;
wire nc30806;
wire nc30807;
wire nc30808;
wire nc30809;
wire nc30810;
wire nc30811;
wire nc30812;
wire nc30813;
wire nc30814;
wire nc30815;
wire nc30816;
wire nc30817;
wire nc30818;
wire nc30819;
wire nc30820;
wire nc30821;
wire nc30822;
wire nc30823;
wire nc30824;
wire nc30825;
wire nc30826;
wire nc30827;
wire nc30828;
wire nc30829;
wire nc30830;
wire nc30831;
wire nc30832;
wire nc30833;
wire nc30834;
wire nc30835;
wire nc30836;
wire nc30837;
wire nc30838;
wire nc30839;
wire nc30840;
wire nc30841;
wire nc30842;
wire nc30843;
wire nc30844;
wire nc30845;
wire nc30846;
wire nc30847;
wire nc30848;
wire nc30849;
wire nc30850;
wire nc30851;
wire nc30852;
wire nc30853;
wire nc30854;
wire nc30855;
wire nc30856;
wire nc30857;
wire nc30858;
wire nc30859;
wire nc30860;
wire nc30861;
wire nc30862;
wire nc30863;
wire nc30864;
wire nc30865;
wire nc30866;
wire nc30867;
wire nc30868;
wire nc30869;
wire nc30870;
wire nc30871;
wire nc30872;
wire nc30873;
wire nc30874;
wire nc30875;
wire nc30876;
wire nc30877;
wire nc30878;
wire nc30879;
wire nc30880;
wire nc30881;
wire nc30882;
wire nc30883;
wire nc30884;
wire nc30885;
wire nc30886;
wire nc30887;
wire nc30888;
wire nc30889;
wire nc30890;
wire nc30891;
wire nc30892;
wire nc30893;
wire nc30894;
wire nc30895;
wire nc30896;
wire nc30897;
wire nc30898;
wire nc30899;
wire nc30900;
wire nc30901;
wire nc30902;
wire nc30903;
wire nc30904;
wire nc30905;
wire nc30906;
wire nc30907;
wire nc30908;
wire nc30909;
wire nc30910;
wire nc30911;
wire nc30912;
wire nc30913;
wire nc30914;
wire nc30915;
wire nc30916;
wire nc30917;
wire nc30918;
wire nc30919;
wire nc30920;
wire nc30921;
wire nc30922;
wire nc30923;
wire nc30924;
wire nc30925;
wire nc30926;
wire nc30927;
wire nc30928;
wire nc30929;
wire nc30930;
wire nc30931;
wire nc30932;
wire nc30933;
wire nc30934;
wire nc30935;
wire nc30936;
wire nc30937;
wire nc30938;
wire nc30939;
wire nc30940;
wire nc30941;
wire nc30942;
wire nc30943;
wire nc30944;
wire nc30945;
wire nc30946;
wire nc30947;
wire nc30948;
wire nc30949;
wire nc30950;
wire nc30951;
wire nc30952;
wire nc30953;
wire nc30954;
wire nc30955;
wire nc30956;
wire nc30957;
wire nc30958;
wire nc30959;
wire nc30960;
wire nc30961;
wire nc30962;
wire nc30963;
wire nc30964;
wire nc30965;
wire nc30966;
wire nc30967;
wire nc30968;
wire nc30969;
wire nc30970;
wire nc30971;
wire nc30972;
wire nc30973;
wire nc30974;
wire nc30975;
wire nc30976;
wire nc30977;
wire nc30978;
wire nc30979;
wire nc30980;
wire nc30981;
wire nc30982;
wire nc30983;
wire nc30984;
wire nc30985;
wire nc30986;
wire nc30987;
wire nc30988;
wire nc30989;
wire nc30990;
wire nc30991;
wire nc30992;
wire nc30993;
wire nc30994;
wire nc30995;
wire nc30996;
wire nc30997;
wire nc30998;
wire nc30999;
wire nc31000;
wire nc31001;
wire nc31002;
wire nc31003;
wire nc31004;
wire nc31005;
wire nc31006;
wire nc31007;
wire nc31008;
wire nc31009;
wire nc31010;
wire nc31011;
wire nc31012;
wire nc31013;
wire nc31014;
wire nc31015;
wire nc31016;
wire nc31017;
wire nc31018;
wire nc31019;
wire nc31020;
wire nc31021;
wire nc31022;
wire nc31023;
wire nc31024;
wire nc31025;
wire nc31026;
wire nc31027;
wire nc31028;
wire nc31029;
wire nc31030;
wire nc31031;
wire nc31032;
wire nc31033;
wire nc31034;
wire nc31035;
wire nc31036;
wire nc31037;
wire nc31038;
wire nc31039;
wire nc31040;
wire nc31041;
wire nc31042;
wire nc31043;
wire nc31044;
wire nc31045;
wire nc31046;
wire nc31047;
wire nc31048;
wire nc31049;
wire nc31050;
wire nc31051;
wire nc31052;
wire nc31053;
wire nc31054;
wire nc31055;
wire nc31056;
wire nc31057;
wire nc31058;
wire nc31059;
wire nc31060;
wire nc31061;
wire nc31062;
wire nc31063;
wire nc31064;
wire nc31065;
wire nc31066;
wire nc31067;
wire nc31068;
wire nc31069;
wire nc31070;
wire nc31071;
wire nc31072;
wire nc31073;
wire nc31074;
wire nc31075;
wire nc31076;
wire nc31077;
wire nc31078;
wire nc31079;
wire nc31080;
wire nc31081;
wire nc31082;
wire nc31083;
wire nc31084;
wire nc31085;
wire nc31086;
wire nc31087;
wire nc31088;
wire nc31089;
wire nc31090;
wire nc31091;
wire nc31092;
wire nc31093;
wire nc31094;
wire nc31095;
wire nc31096;
wire nc31097;
wire nc31098;
wire nc31099;
wire nc31100;
wire nc31101;
wire nc31102;
wire nc31103;
wire nc31104;
wire nc31105;
wire nc31106;
wire nc31107;
wire nc31108;
wire nc31109;
wire nc31110;
wire nc31111;
wire nc31112;
wire nc31113;
wire nc31114;
wire nc31115;
wire nc31116;
wire nc31117;
wire nc31118;
wire nc31119;
wire nc31120;
wire nc31121;
wire nc31122;
wire nc31123;
wire nc31124;
wire nc31125;
wire nc31126;
wire nc31127;
wire nc31128;
wire nc31129;
wire nc31130;
wire nc31131;
wire nc31132;
wire nc31133;
wire nc31134;
wire nc31135;
wire nc31136;
wire nc31137;
wire nc31138;
wire nc31139;
wire nc31140;
wire nc31141;
wire nc31142;
wire nc31143;
wire nc31144;
wire nc31145;
wire nc31146;
wire nc31147;
wire nc31148;
wire nc31149;
wire nc31150;
wire nc31151;
wire nc31152;
wire nc31153;
wire nc31154;
wire nc31155;
wire nc31156;
wire nc31157;
wire nc31158;
wire nc31159;
wire nc31160;
wire nc31161;
wire nc31162;
wire nc31163;
wire nc31164;
wire nc31165;
wire nc31166;
wire nc31167;
wire nc31168;
wire nc31169;
wire nc31170;
wire nc31171;
wire nc31172;
wire nc31173;
wire nc31174;
wire nc31175;
wire nc31176;
wire nc31177;
wire nc31178;
wire nc31179;
wire nc31180;
wire nc31181;
wire nc31182;
wire nc31183;
wire nc31184;
wire nc31185;
wire nc31186;
wire nc31187;
wire nc31188;
wire nc31189;
wire nc31190;
wire nc31191;
wire nc31192;
wire nc31193;
wire nc31194;
wire nc31195;
wire nc31196;
wire nc31197;
wire nc31198;
wire nc31199;
wire nc31200;
wire nc31201;
wire nc31202;
wire nc31203;
wire nc31204;
wire nc31205;
wire nc31206;
wire nc31207;
wire nc31208;
wire nc31209;
wire nc31210;
wire nc31211;
wire nc31212;
wire nc31213;
wire nc31214;
wire nc31215;
wire nc31216;
wire nc31217;
wire nc31218;
wire nc31219;
wire nc31220;
wire nc31221;
wire nc31222;
wire nc31223;
wire nc31224;
wire nc31225;
wire nc31226;
wire nc31227;
wire nc31228;
wire nc31229;
wire nc31230;
wire nc31231;
wire nc31232;
wire nc31233;
wire nc31234;
wire nc31235;
wire nc31236;
wire nc31237;
wire nc31238;
wire nc31239;
wire nc31240;
wire nc31241;
wire nc31242;
wire nc31243;
wire nc31244;
wire nc31245;
wire nc31246;
wire nc31247;
wire nc31248;
wire nc31249;
wire nc31250;
wire nc31251;
wire nc31252;
wire nc31253;
wire nc31254;
wire nc31255;
wire nc31256;
wire nc31257;
wire nc31258;
wire nc31259;
wire nc31260;
wire nc31261;
wire nc31262;
wire nc31263;
wire nc31264;
wire nc31265;
wire nc31266;
wire nc31267;
wire nc31268;
wire nc31269;
wire nc31270;
wire nc31271;
wire nc31272;
wire nc31273;
wire nc31274;
wire nc31275;
wire nc31276;
wire nc31277;
wire nc31278;
wire nc31279;
wire nc31280;
wire nc31281;
wire nc31282;
wire nc31283;
wire nc31284;
wire nc31285;
wire nc31286;
wire nc31287;
wire nc31288;
wire nc31289;
wire nc31290;
wire nc31291;
wire nc31292;
wire nc31293;
wire nc31294;
wire nc31295;
wire nc31296;
wire nc31297;
wire nc31298;
wire nc31299;
wire nc31300;
wire nc31301;
wire nc31302;
wire nc31303;
wire nc31304;
wire nc31305;
wire nc31306;
wire nc31307;
wire nc31308;
wire nc31309;
wire nc31310;
wire nc31311;
wire nc31312;
wire nc31313;
wire nc31314;
wire nc31315;
wire nc31316;
wire nc31317;
wire nc31318;
wire nc31319;
wire nc31320;
wire nc31321;
wire nc31322;
wire nc31323;
wire nc31324;
wire nc31325;
wire nc31326;
wire nc31327;
wire nc31328;
wire nc31329;
wire nc31330;
wire nc31331;
wire nc31332;
wire nc31333;
wire nc31334;
wire nc31335;
wire nc31336;
wire nc31337;
wire nc31338;
wire nc31339;
wire nc31340;
wire nc31341;
wire nc31342;
wire nc31343;
wire nc31344;
wire nc31345;
wire nc31346;
wire nc31347;
wire nc31348;
wire nc31349;
wire nc31350;
wire nc31351;
wire nc31352;
wire nc31353;
wire nc31354;
wire nc31355;
wire nc31356;
wire nc31357;
wire nc31358;
wire nc31359;
wire nc31360;
wire nc31361;
wire nc31362;
wire nc31363;
wire nc31364;
wire nc31365;
wire nc31366;
wire nc31367;
wire nc31368;
wire nc31369;
wire nc31370;
wire nc31371;
wire nc31372;
wire nc31373;
wire nc31374;
wire nc31375;
wire nc31376;
wire nc31377;
wire nc31378;
wire nc31379;
wire nc31380;
wire nc31381;
wire nc31382;
wire nc31383;
wire nc31384;
wire nc31385;
wire nc31386;
wire nc31387;
wire nc31388;
wire nc31389;
wire nc31390;
wire nc31391;
wire nc31392;
wire nc31393;
wire nc31394;
wire nc31395;
wire nc31396;
wire nc31397;
wire nc31398;
wire nc31399;
wire nc31400;
wire nc31401;
wire nc31402;
wire nc31403;
wire nc31404;
wire nc31405;
wire nc31406;
wire nc31407;
wire nc31408;
wire nc31409;
wire nc31410;
wire nc31411;
wire nc31412;
wire nc31413;
wire nc31414;
wire nc31415;
wire nc31416;
wire nc31417;
wire nc31418;
wire nc31419;
wire nc31420;
wire nc31421;
wire nc31422;
wire nc31423;
wire nc31424;
wire nc31425;
wire nc31426;
wire nc31427;
wire nc31428;
wire nc31429;
wire nc31430;
wire nc31431;
wire nc31432;
wire nc31433;
wire nc31434;
wire nc31435;
wire nc31436;
wire nc31437;
wire nc31438;
wire nc31439;
wire nc31440;
wire nc31441;
wire nc31442;
wire nc31443;
wire nc31444;
wire nc31445;
wire nc31446;
wire nc31447;
wire nc31448;
wire nc31449;
wire nc31450;
wire nc31451;
wire nc31452;
wire nc31453;
wire nc31454;
wire nc31455;
wire nc31456;
wire nc31457;
wire nc31458;
wire nc31459;
wire nc31460;
wire nc31461;
wire nc31462;
wire nc31463;
wire nc31464;
wire nc31465;
wire nc31466;
wire nc31467;
wire nc31468;
wire nc31469;
wire nc31470;
wire nc31471;
wire nc31472;
wire nc31473;
wire nc31474;
wire nc31475;
wire nc31476;
wire nc31477;
wire nc31478;
wire nc31479;
wire nc31480;
wire nc31481;
wire nc31482;
wire nc31483;
wire nc31484;
wire nc31485;
wire nc31486;
wire nc31487;
wire nc31488;
wire nc31489;
wire nc31490;
wire nc31491;
wire nc31492;
wire nc31493;
wire nc31494;
wire nc31495;
wire nc31496;
wire nc31497;
wire nc31498;
wire nc31499;
wire nc31500;
wire nc31501;
wire nc31502;
wire nc31503;
wire nc31504;
wire nc31505;
wire nc31506;
wire nc31507;
wire nc31508;
wire nc31509;
wire nc31510;
wire nc31511;
wire nc31512;
wire nc31513;
wire nc31514;
wire nc31515;
wire nc31516;
wire nc31517;
wire nc31518;
wire nc31519;
wire nc31520;
wire nc31521;
wire nc31522;
wire nc31523;
wire nc31524;
wire nc31525;
wire nc31526;
wire nc31527;
wire nc31528;
wire nc31529;
wire nc31530;
wire nc31531;
wire nc31532;
wire nc31533;
wire nc31534;
wire nc31535;
wire nc31536;
wire nc31537;
wire nc31538;
wire nc31539;
wire nc31540;
wire nc31541;
wire nc31542;
wire nc31543;
wire nc31544;
wire nc31545;
wire nc31546;
wire nc31547;
wire nc31548;
wire nc31549;
wire nc31550;
wire nc31551;
wire nc31552;
wire nc31553;
wire nc31554;
wire nc31555;
wire nc31556;
wire nc31557;
wire nc31558;
wire nc31559;
wire nc31560;
wire nc31561;
wire nc31562;
wire nc31563;
wire nc31564;
wire nc31565;
wire nc31566;
wire nc31567;
wire nc31568;
wire nc31569;
wire nc31570;
wire nc31571;
wire nc31572;
wire nc31573;
wire nc31574;
wire nc31575;
wire nc31576;
wire nc31577;
wire nc31578;
wire nc31579;
wire nc31580;
wire nc31581;
wire nc31582;
wire nc31583;
wire nc31584;
wire nc31585;
wire nc31586;
wire nc31587;
wire nc31588;
wire nc31589;
wire nc31590;
wire nc31591;
wire nc31592;
wire nc31593;
wire nc31594;
wire nc31595;
wire nc31596;
wire nc31597;
wire nc31598;
wire nc31599;
wire nc31600;
wire nc31601;
wire nc31602;
wire nc31603;
wire nc31604;
wire nc31605;
wire nc31606;
wire nc31607;
wire nc31608;
wire nc31609;
wire nc31610;
wire nc31611;
wire nc31612;
wire nc31613;
wire nc31614;
wire nc31615;
wire nc31616;
wire nc31617;
wire nc31618;
wire nc31619;
wire nc31620;
wire nc31621;
wire nc31622;
wire nc31623;
wire nc31624;
wire nc31625;
wire nc31626;
wire nc31627;
wire nc31628;
wire nc31629;
wire nc31630;
wire nc31631;
wire nc31632;
wire nc31633;
wire nc31634;
wire nc31635;
wire nc31636;
wire nc31637;
wire nc31638;
wire nc31639;
wire nc31640;
wire nc31641;
wire nc31642;
wire nc31643;
wire nc31644;
wire nc31645;
wire nc31646;
wire nc31647;
wire nc31648;
wire nc31649;
wire nc31650;
wire nc31651;
wire nc31652;
wire nc31653;
wire nc31654;
wire nc31655;
wire nc31656;
wire nc31657;
wire nc31658;
wire nc31659;
wire nc31660;
wire nc31661;
wire nc31662;
wire nc31663;
wire nc31664;
wire nc31665;
wire nc31666;
wire nc31667;
wire nc31668;
wire nc31669;
wire nc31670;
wire nc31671;
wire nc31672;
wire nc31673;
wire nc31674;
wire nc31675;
wire nc31676;
wire nc31677;
wire nc31678;
wire nc31679;
wire nc31680;
wire nc31681;
wire nc31682;
wire nc31683;
wire nc31684;
wire nc31685;
wire nc31686;
wire nc31687;
wire nc31688;
wire nc31689;
wire nc31690;
wire nc31691;
wire nc31692;
wire nc31693;
wire nc31694;
wire nc31695;
wire nc31696;
wire nc31697;
wire nc31698;
wire nc31699;
wire nc31700;
wire nc31701;
wire nc31702;
wire nc31703;
wire nc31704;
wire nc31705;
wire nc31706;
wire nc31707;
wire nc31708;
wire nc31709;
wire nc31710;
wire nc31711;
wire nc31712;
wire nc31713;
wire nc31714;
wire nc31715;
wire nc31716;
wire nc31717;
wire nc31718;
wire nc31719;
wire nc31720;
wire nc31721;
wire nc31722;
wire nc31723;
wire nc31724;
wire nc31725;
wire nc31726;
wire nc31727;
wire nc31728;
wire nc31729;
wire nc31730;
wire nc31731;
wire nc31732;
wire nc31733;
wire nc31734;
wire nc31735;
wire nc31736;
wire nc31737;
wire nc31738;
wire nc31739;
wire nc31740;
wire nc31741;
wire nc31742;
wire nc31743;
wire nc31744;
wire nc31745;
wire nc31746;
wire nc31747;
wire nc31748;
wire nc31749;
wire nc31750;
wire nc31751;
wire nc31752;
wire nc31753;
wire nc31754;
wire nc31755;
wire nc31756;
wire nc31757;
wire nc31758;
wire nc31759;
wire nc31760;
wire nc31761;
wire nc31762;
wire nc31763;
wire nc31764;
wire nc31765;
wire nc31766;
wire nc31767;
wire nc31768;
wire nc31769;
wire nc31770;
wire nc31771;
wire nc31772;
wire nc31773;
wire nc31774;
wire nc31775;
wire nc31776;
wire nc31777;
wire nc31778;
wire nc31779;
wire nc31780;
wire nc31781;
wire nc31782;
wire nc31783;
wire nc31784;
wire nc31785;
wire nc31786;
wire nc31787;
wire nc31788;
wire nc31789;
wire nc31790;
wire nc31791;
wire nc31792;
wire nc31793;
wire nc31794;
wire nc31795;
wire nc31796;
wire nc31797;
wire nc31798;
wire nc31799;
wire nc31800;
wire nc31801;
wire nc31802;
wire nc31803;
wire nc31804;
wire nc31805;
wire nc31806;
wire nc31807;
wire nc31808;
wire nc31809;
wire nc31810;
wire nc31811;
wire nc31812;
wire nc31813;
wire nc31814;
wire nc31815;
wire nc31816;
wire nc31817;
wire nc31818;
wire nc31819;
wire nc31820;
wire nc31821;
wire nc31822;
wire nc31823;
wire nc31824;
wire nc31825;
wire nc31826;
wire nc31827;
wire nc31828;
wire nc31829;
wire nc31830;
wire nc31831;
wire nc31832;
wire nc31833;
wire nc31834;
wire nc31835;
wire nc31836;
wire nc31837;
wire nc31838;
wire nc31839;
wire nc31840;
wire nc31841;
wire nc31842;
wire nc31843;
wire nc31844;
wire nc31845;
wire nc31846;
wire nc31847;
wire nc31848;
wire nc31849;
wire nc31850;
wire nc31851;
wire nc31852;
wire nc31853;
wire nc31854;
wire nc31855;
wire nc31856;
wire nc31857;
wire nc31858;
wire nc31859;
wire nc31860;
wire nc31861;
wire nc31862;
wire nc31863;
wire nc31864;
wire nc31865;
wire nc31866;
wire nc31867;
wire nc31868;
wire nc31869;
wire nc31870;
wire nc31871;
wire nc31872;
wire nc31873;
wire nc31874;
wire nc31875;
wire nc31876;
wire nc31877;
wire nc31878;
wire nc31879;
wire nc31880;
wire nc31881;
wire nc31882;
wire nc31883;
wire nc31884;
wire nc31885;
wire nc31886;
wire nc31887;
wire nc31888;
wire nc31889;
wire nc31890;
wire nc31891;
wire nc31892;
wire nc31893;
wire nc31894;
wire nc31895;
wire nc31896;
wire nc31897;
wire nc31898;
wire nc31899;
wire nc31900;
wire nc31901;
wire nc31902;
wire nc31903;
wire nc31904;
wire nc31905;
wire nc31906;
wire nc31907;
wire nc31908;
wire nc31909;
wire nc31910;
wire nc31911;
wire nc31912;
wire nc31913;
wire nc31914;
wire nc31915;
wire nc31916;
wire nc31917;
wire nc31918;
wire nc31919;
wire nc31920;
wire nc31921;
wire nc31922;
wire nc31923;
wire nc31924;
wire nc31925;
wire nc31926;
wire nc31927;
wire nc31928;
wire nc31929;
wire nc31930;
wire nc31931;
wire nc31932;
wire nc31933;
wire nc31934;
wire nc31935;
wire nc31936;
wire nc31937;
wire nc31938;
wire nc31939;
wire nc31940;
wire nc31941;
wire nc31942;
wire nc31943;
wire nc31944;
wire nc31945;
wire nc31946;
wire nc31947;
wire nc31948;
wire nc31949;
wire nc31950;
wire nc31951;
wire nc31952;
wire nc31953;
wire nc31954;
wire nc31955;
wire nc31956;
wire nc31957;
wire nc31958;
wire nc31959;
wire nc31960;
wire nc31961;
wire nc31962;
wire nc31963;
wire nc31964;
wire nc31965;
wire nc31966;
wire nc31967;
wire nc31968;
wire nc31969;
wire nc31970;
wire nc31971;
wire nc31972;
wire nc31973;
wire nc31974;
wire nc31975;
wire nc31976;
wire nc31977;
wire nc31978;
wire nc31979;
wire nc31980;
wire nc31981;
wire nc31982;
wire nc31983;
wire nc31984;
wire nc31985;
wire nc31986;
wire nc31987;
wire nc31988;
wire nc31989;
wire nc31990;
wire nc31991;
wire nc31992;
wire nc31993;
wire nc31994;
wire nc31995;
wire nc31996;
wire nc31997;
wire nc31998;
wire nc31999;
wire nc32000;
wire nc32001;
wire nc32002;
wire nc32003;
wire nc32004;
wire nc32005;
wire nc32006;
wire nc32007;
wire nc32008;
wire nc32009;
wire nc32010;
wire nc32011;
wire nc32012;
wire nc32013;
wire nc32014;
wire nc32015;
wire nc32016;
wire nc32017;
wire nc32018;
wire nc32019;
wire nc32020;
wire nc32021;
wire nc32022;
wire nc32023;
wire nc32024;
wire nc32025;
wire nc32026;
wire nc32027;
wire nc32028;
wire nc32029;
wire nc32030;
wire nc32031;
wire nc32032;
wire nc32033;
wire nc32034;
wire nc32035;
wire nc32036;
wire nc32037;
wire nc32038;
wire nc32039;
wire nc32040;
wire nc32041;
wire nc32042;
wire nc32043;
wire nc32044;
wire nc32045;
wire nc32046;
wire nc32047;
wire nc32048;
wire nc32049;
wire nc32050;
wire nc32051;
wire nc32052;
wire nc32053;
wire nc32054;
wire nc32055;
wire nc32056;
wire nc32057;
wire nc32058;
wire nc32059;
wire nc32060;
wire nc32061;
wire nc32062;
wire nc32063;
wire nc32064;
wire nc32065;
wire nc32066;
wire nc32067;
wire nc32068;
wire nc32069;
wire nc32070;
wire nc32071;
wire nc32072;
wire nc32073;
wire nc32074;
wire nc32075;
wire nc32076;
wire nc32077;
wire nc32078;
wire nc32079;
wire nc32080;
wire nc32081;
wire nc32082;
wire nc32083;
wire nc32084;
wire nc32085;
wire nc32086;
wire nc32087;
wire nc32088;
wire nc32089;
wire nc32090;
wire nc32091;
wire nc32092;
wire nc32093;
wire nc32094;
wire nc32095;
wire nc32096;
wire nc32097;
wire nc32098;
wire nc32099;
wire nc32100;
wire nc32101;
wire nc32102;
wire nc32103;
wire nc32104;
wire nc32105;
wire nc32106;
wire nc32107;
wire nc32108;
wire nc32109;
wire nc32110;
wire nc32111;
wire nc32112;
wire nc32113;
wire nc32114;
wire nc32115;
wire nc32116;
wire nc32117;
wire nc32118;
wire nc32119;
wire nc32120;
wire nc32121;
wire nc32122;
wire nc32123;
wire nc32124;
wire nc32125;
wire nc32126;
wire nc32127;
wire nc32128;
wire nc32129;
wire nc32130;
wire nc32131;
wire nc32132;
wire nc32133;
wire nc32134;
wire nc32135;
wire nc32136;
wire nc32137;
wire nc32138;
wire nc32139;
wire nc32140;
wire nc32141;
wire nc32142;
wire nc32143;
wire nc32144;
wire nc32145;
wire nc32146;
wire nc32147;
wire nc32148;
wire nc32149;
wire nc32150;
wire nc32151;
wire nc32152;
wire nc32153;
wire nc32154;
wire nc32155;
wire nc32156;
wire nc32157;
wire nc32158;
wire nc32159;
wire nc32160;
wire nc32161;
wire nc32162;
wire nc32163;
wire nc32164;
wire nc32165;
wire nc32166;
wire nc32167;
wire nc32168;
wire nc32169;
wire nc32170;
wire nc32171;
wire nc32172;
wire nc32173;
wire nc32174;
wire nc32175;
wire nc32176;
wire nc32177;
wire nc32178;
wire nc32179;
wire nc32180;
wire nc32181;
wire nc32182;
wire nc32183;
wire nc32184;
wire nc32185;
wire nc32186;
wire nc32187;
wire nc32188;
wire nc32189;
wire nc32190;
wire nc32191;
wire nc32192;
wire nc32193;
wire nc32194;
wire nc32195;
wire nc32196;
wire nc32197;
wire nc32198;
wire nc32199;
wire nc32200;
wire nc32201;
wire nc32202;
wire nc32203;
wire nc32204;
wire nc32205;
wire nc32206;
wire nc32207;
wire nc32208;
wire nc32209;
wire nc32210;
wire nc32211;
wire nc32212;
wire nc32213;
wire nc32214;
wire nc32215;
wire nc32216;
wire nc32217;
wire nc32218;
wire nc32219;
wire nc32220;
wire nc32221;
wire nc32222;
wire nc32223;
wire nc32224;
wire nc32225;
wire nc32226;
wire nc32227;
wire nc32228;
wire nc32229;
wire nc32230;
wire nc32231;
wire nc32232;
wire nc32233;
wire nc32234;
wire nc32235;
wire nc32236;
wire nc32237;
wire nc32238;
wire nc32239;
wire nc32240;
wire nc32241;
wire nc32242;
wire nc32243;
wire nc32244;
wire nc32245;
wire nc32246;
wire nc32247;
wire nc32248;
wire nc32249;
wire nc32250;
wire nc32251;
wire nc32252;
wire nc32253;
wire nc32254;
wire nc32255;
wire nc32256;

assign vcc_net = 1;
assign gnd_net = 0;
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_0 (
		.doa ({nc16129, nc16130, nc16131, nc16132, nc16133, nc16134, nc16135, nc16136, nc16137, nc16138, nc16139, nc16140, nc16141, nc16142, nc16143, nc16144, nc16145, nc16146, nc16147, nc16148, nc16149, nc16150, nc16151, nc16152, nc16153, nc16154, nc16155, nc16156, nc16157, nc16158, nc16159, nc16160, nc16161, nc16162, nc16163, nc16164, nc16165, nc16166, nc16167, nc16168, nc16169, nc16170, nc16171, nc16172, nc16173, nc16174, nc16175, nc16176, nc16177, nc16178, nc16179, nc16180, nc16181, nc16182, nc16183, nc16184, nc16185, nc16186, nc16187, nc16188, nc16189, nc16190, nc16191, net_33}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc16192, nc16193, nc16194, nc16195, nc16196, nc16197, nc16198, nc16199, nc16200, nc16201, nc16202, nc16203, nc16204, nc16205, nc16206, nc16207, nc16208, nc16209, nc16210, nc16211, nc16212, nc16213, nc16214, nc16215, nc16216, nc16217, nc16218, nc16219, nc16220, nc16221, nc16222, nc16223, nc16224, nc16225, nc16226, nc16227, nc16228, nc16229, nc16230, nc16231, nc16232, nc16233, nc16234, nc16235, nc16236, nc16237, nc16238, nc16239, nc16240, nc16241, nc16242, nc16243, nc16244, nc16245, nc16246, nc16247, nc16248, nc16249, nc16250, nc16251, nc16252, nc16253, nc16254, dw[0]}),
		.dipa (),
		.dipb (),
		.cea (net_3),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_4 (
		.doa ({nc16255, nc16256, nc16257, nc16258, nc16259, nc16260, nc16261, nc16262, nc16263, nc16264, nc16265, nc16266, nc16267, nc16268, nc16269, nc16270, nc16271, nc16272, nc16273, nc16274, nc16275, nc16276, nc16277, nc16278, nc16279, nc16280, nc16281, nc16282, nc16283, nc16284, nc16285, nc16286, nc16287, nc16288, nc16289, nc16290, nc16291, nc16292, nc16293, nc16294, nc16295, nc16296, nc16297, nc16298, nc16299, nc16300, nc16301, nc16302, nc16303, nc16304, nc16305, nc16306, nc16307, nc16308, nc16309, nc16310, nc16311, nc16312, nc16313, nc16314, nc16315, nc16316, nc16317, net_37}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc16318, nc16319, nc16320, nc16321, nc16322, nc16323, nc16324, nc16325, nc16326, nc16327, nc16328, nc16329, nc16330, nc16331, nc16332, nc16333, nc16334, nc16335, nc16336, nc16337, nc16338, nc16339, nc16340, nc16341, nc16342, nc16343, nc16344, nc16345, nc16346, nc16347, nc16348, nc16349, nc16350, nc16351, nc16352, nc16353, nc16354, nc16355, nc16356, nc16357, nc16358, nc16359, nc16360, nc16361, nc16362, nc16363, nc16364, nc16365, nc16366, nc16367, nc16368, nc16369, nc16370, nc16371, nc16372, nc16373, nc16374, nc16375, nc16376, nc16377, nc16378, nc16379, nc16380, dw[8]}),
		.dipa (),
		.dipb (),
		.cea (net_35),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_ADDR_PIPE_A u_addra_pipe_0 (
		.clk (clkr),
		.ena (cer),
		.i (ar[0]),
		.o (addra_pipe_0_net)
	);
fifo2ram_emb_v1_MUX u0 (
		.sel (addra_pipe_0_net),
		.i0 (net_33),
		.i1 (net_37),
		.o (net_41)
	);
fifo2ram_emb_v1_AND u1 (
		.i0 (net_43),
		.i1 (net_42),
		.o (net_3)
	);
fifo2ram_emb_v1_AND u2 (
		.i0 (net_43),
		.i1 (ar[0]),
		.o (net_35)
	);
fifo2ram_emb_v1_NOT u3 (
		.i (ar[0]),
		.o (net_42)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_8 (
		.doa ({nc16381, nc16382, nc16383, nc16384, nc16385, nc16386, nc16387, nc16388, nc16389, nc16390, nc16391, nc16392, nc16393, nc16394, nc16395, nc16396, nc16397, nc16398, nc16399, nc16400, nc16401, nc16402, nc16403, nc16404, nc16405, nc16406, nc16407, nc16408, nc16409, nc16410, nc16411, nc16412, nc16413, nc16414, nc16415, nc16416, nc16417, nc16418, nc16419, nc16420, nc16421, nc16422, nc16423, nc16424, nc16425, nc16426, nc16427, nc16428, nc16429, nc16430, nc16431, nc16432, nc16433, nc16434, nc16435, nc16436, nc16437, nc16438, nc16439, nc16440, nc16441, nc16442, nc16443, net_46}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc16444, nc16445, nc16446, nc16447, nc16448, nc16449, nc16450, nc16451, nc16452, nc16453, nc16454, nc16455, nc16456, nc16457, nc16458, nc16459, nc16460, nc16461, nc16462, nc16463, nc16464, nc16465, nc16466, nc16467, nc16468, nc16469, nc16470, nc16471, nc16472, nc16473, nc16474, nc16475, nc16476, nc16477, nc16478, nc16479, nc16480, nc16481, nc16482, nc16483, nc16484, nc16485, nc16486, nc16487, nc16488, nc16489, nc16490, nc16491, nc16492, nc16493, nc16494, nc16495, nc16496, nc16497, nc16498, nc16499, nc16500, nc16501, nc16502, nc16503, nc16504, nc16505, nc16506, dw[16]}),
		.dipa (),
		.dipb (),
		.cea (net_44),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_12 (
		.doa ({nc16507, nc16508, nc16509, nc16510, nc16511, nc16512, nc16513, nc16514, nc16515, nc16516, nc16517, nc16518, nc16519, nc16520, nc16521, nc16522, nc16523, nc16524, nc16525, nc16526, nc16527, nc16528, nc16529, nc16530, nc16531, nc16532, nc16533, nc16534, nc16535, nc16536, nc16537, nc16538, nc16539, nc16540, nc16541, nc16542, nc16543, nc16544, nc16545, nc16546, nc16547, nc16548, nc16549, nc16550, nc16551, nc16552, nc16553, nc16554, nc16555, nc16556, nc16557, nc16558, nc16559, nc16560, nc16561, nc16562, nc16563, nc16564, nc16565, nc16566, nc16567, nc16568, nc16569, net_50}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc16570, nc16571, nc16572, nc16573, nc16574, nc16575, nc16576, nc16577, nc16578, nc16579, nc16580, nc16581, nc16582, nc16583, nc16584, nc16585, nc16586, nc16587, nc16588, nc16589, nc16590, nc16591, nc16592, nc16593, nc16594, nc16595, nc16596, nc16597, nc16598, nc16599, nc16600, nc16601, nc16602, nc16603, nc16604, nc16605, nc16606, nc16607, nc16608, nc16609, nc16610, nc16611, nc16612, nc16613, nc16614, nc16615, nc16616, nc16617, nc16618, nc16619, nc16620, nc16621, nc16622, nc16623, nc16624, nc16625, nc16626, nc16627, nc16628, nc16629, nc16630, nc16631, nc16632, dw[24]}),
		.dipa (),
		.dipb (),
		.cea (net_48),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u4 (
		.sel (addra_pipe_0_net),
		.i0 (net_46),
		.i1 (net_50),
		.o (net_52)
	);
fifo2ram_emb_v1_AND u5 (
		.i0 (net_54),
		.i1 (net_53),
		.o (net_44)
	);
fifo2ram_emb_v1_AND u6 (
		.i0 (net_54),
		.i1 (ar[0]),
		.o (net_48)
	);
fifo2ram_emb_v1_NOT u7 (
		.i (ar[0]),
		.o (net_53)
	);
fifo2ram_emb_v1_ADDR_PIPE_A u_addra_pipe_1 (
		.clk (clkr),
		.ena (cer),
		.i (ar[1]),
		.o (addra_pipe_1_net)
	);
fifo2ram_emb_v1_MUX u8 (
		.sel (addra_pipe_1_net),
		.i0 (net_41),
		.i1 (net_52),
		.o (net_56)
	);
fifo2ram_emb_v1_AND u9 (
		.i0 (net_58),
		.i1 (net_57),
		.o (net_43)
	);
fifo2ram_emb_v1_AND u10 (
		.i0 (net_58),
		.i1 (ar[1]),
		.o (net_54)
	);
fifo2ram_emb_v1_NOT u11 (
		.i (ar[1]),
		.o (net_57)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_16 (
		.doa ({nc16633, nc16634, nc16635, nc16636, nc16637, nc16638, nc16639, nc16640, nc16641, nc16642, nc16643, nc16644, nc16645, nc16646, nc16647, nc16648, nc16649, nc16650, nc16651, nc16652, nc16653, nc16654, nc16655, nc16656, nc16657, nc16658, nc16659, nc16660, nc16661, nc16662, nc16663, nc16664, nc16665, nc16666, nc16667, nc16668, nc16669, nc16670, nc16671, nc16672, nc16673, nc16674, nc16675, nc16676, nc16677, nc16678, nc16679, nc16680, nc16681, nc16682, nc16683, nc16684, nc16685, nc16686, nc16687, nc16688, nc16689, nc16690, nc16691, nc16692, nc16693, nc16694, nc16695, net_61}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc16696, nc16697, nc16698, nc16699, nc16700, nc16701, nc16702, nc16703, nc16704, nc16705, nc16706, nc16707, nc16708, nc16709, nc16710, nc16711, nc16712, nc16713, nc16714, nc16715, nc16716, nc16717, nc16718, nc16719, nc16720, nc16721, nc16722, nc16723, nc16724, nc16725, nc16726, nc16727, nc16728, nc16729, nc16730, nc16731, nc16732, nc16733, nc16734, nc16735, nc16736, nc16737, nc16738, nc16739, nc16740, nc16741, nc16742, nc16743, nc16744, nc16745, nc16746, nc16747, nc16748, nc16749, nc16750, nc16751, nc16752, nc16753, nc16754, nc16755, nc16756, nc16757, nc16758, dw[32]}),
		.dipa (),
		.dipb (),
		.cea (net_59),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_20 (
		.doa ({nc16759, nc16760, nc16761, nc16762, nc16763, nc16764, nc16765, nc16766, nc16767, nc16768, nc16769, nc16770, nc16771, nc16772, nc16773, nc16774, nc16775, nc16776, nc16777, nc16778, nc16779, nc16780, nc16781, nc16782, nc16783, nc16784, nc16785, nc16786, nc16787, nc16788, nc16789, nc16790, nc16791, nc16792, nc16793, nc16794, nc16795, nc16796, nc16797, nc16798, nc16799, nc16800, nc16801, nc16802, nc16803, nc16804, nc16805, nc16806, nc16807, nc16808, nc16809, nc16810, nc16811, nc16812, nc16813, nc16814, nc16815, nc16816, nc16817, nc16818, nc16819, nc16820, nc16821, net_65}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc16822, nc16823, nc16824, nc16825, nc16826, nc16827, nc16828, nc16829, nc16830, nc16831, nc16832, nc16833, nc16834, nc16835, nc16836, nc16837, nc16838, nc16839, nc16840, nc16841, nc16842, nc16843, nc16844, nc16845, nc16846, nc16847, nc16848, nc16849, nc16850, nc16851, nc16852, nc16853, nc16854, nc16855, nc16856, nc16857, nc16858, nc16859, nc16860, nc16861, nc16862, nc16863, nc16864, nc16865, nc16866, nc16867, nc16868, nc16869, nc16870, nc16871, nc16872, nc16873, nc16874, nc16875, nc16876, nc16877, nc16878, nc16879, nc16880, nc16881, nc16882, nc16883, nc16884, dw[40]}),
		.dipa (),
		.dipb (),
		.cea (net_63),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u12 (
		.sel (addra_pipe_0_net),
		.i0 (net_61),
		.i1 (net_65),
		.o (net_67)
	);
fifo2ram_emb_v1_AND u13 (
		.i0 (net_69),
		.i1 (net_68),
		.o (net_59)
	);
fifo2ram_emb_v1_AND u14 (
		.i0 (net_69),
		.i1 (ar[0]),
		.o (net_63)
	);
fifo2ram_emb_v1_NOT u15 (
		.i (ar[0]),
		.o (net_68)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_24 (
		.doa ({nc16885, nc16886, nc16887, nc16888, nc16889, nc16890, nc16891, nc16892, nc16893, nc16894, nc16895, nc16896, nc16897, nc16898, nc16899, nc16900, nc16901, nc16902, nc16903, nc16904, nc16905, nc16906, nc16907, nc16908, nc16909, nc16910, nc16911, nc16912, nc16913, nc16914, nc16915, nc16916, nc16917, nc16918, nc16919, nc16920, nc16921, nc16922, nc16923, nc16924, nc16925, nc16926, nc16927, nc16928, nc16929, nc16930, nc16931, nc16932, nc16933, nc16934, nc16935, nc16936, nc16937, nc16938, nc16939, nc16940, nc16941, nc16942, nc16943, nc16944, nc16945, nc16946, nc16947, net_72}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc16948, nc16949, nc16950, nc16951, nc16952, nc16953, nc16954, nc16955, nc16956, nc16957, nc16958, nc16959, nc16960, nc16961, nc16962, nc16963, nc16964, nc16965, nc16966, nc16967, nc16968, nc16969, nc16970, nc16971, nc16972, nc16973, nc16974, nc16975, nc16976, nc16977, nc16978, nc16979, nc16980, nc16981, nc16982, nc16983, nc16984, nc16985, nc16986, nc16987, nc16988, nc16989, nc16990, nc16991, nc16992, nc16993, nc16994, nc16995, nc16996, nc16997, nc16998, nc16999, nc17000, nc17001, nc17002, nc17003, nc17004, nc17005, nc17006, nc17007, nc17008, nc17009, nc17010, dw[48]}),
		.dipa (),
		.dipb (),
		.cea (net_70),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_28 (
		.doa ({nc17011, nc17012, nc17013, nc17014, nc17015, nc17016, nc17017, nc17018, nc17019, nc17020, nc17021, nc17022, nc17023, nc17024, nc17025, nc17026, nc17027, nc17028, nc17029, nc17030, nc17031, nc17032, nc17033, nc17034, nc17035, nc17036, nc17037, nc17038, nc17039, nc17040, nc17041, nc17042, nc17043, nc17044, nc17045, nc17046, nc17047, nc17048, nc17049, nc17050, nc17051, nc17052, nc17053, nc17054, nc17055, nc17056, nc17057, nc17058, nc17059, nc17060, nc17061, nc17062, nc17063, nc17064, nc17065, nc17066, nc17067, nc17068, nc17069, nc17070, nc17071, nc17072, nc17073, net_76}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17074, nc17075, nc17076, nc17077, nc17078, nc17079, nc17080, nc17081, nc17082, nc17083, nc17084, nc17085, nc17086, nc17087, nc17088, nc17089, nc17090, nc17091, nc17092, nc17093, nc17094, nc17095, nc17096, nc17097, nc17098, nc17099, nc17100, nc17101, nc17102, nc17103, nc17104, nc17105, nc17106, nc17107, nc17108, nc17109, nc17110, nc17111, nc17112, nc17113, nc17114, nc17115, nc17116, nc17117, nc17118, nc17119, nc17120, nc17121, nc17122, nc17123, nc17124, nc17125, nc17126, nc17127, nc17128, nc17129, nc17130, nc17131, nc17132, nc17133, nc17134, nc17135, nc17136, dw[56]}),
		.dipa (),
		.dipb (),
		.cea (net_74),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u16 (
		.sel (addra_pipe_0_net),
		.i0 (net_72),
		.i1 (net_76),
		.o (net_78)
	);
fifo2ram_emb_v1_AND u17 (
		.i0 (net_80),
		.i1 (net_79),
		.o (net_70)
	);
fifo2ram_emb_v1_AND u18 (
		.i0 (net_80),
		.i1 (ar[0]),
		.o (net_74)
	);
fifo2ram_emb_v1_NOT u19 (
		.i (ar[0]),
		.o (net_79)
	);
fifo2ram_emb_v1_MUX u20 (
		.sel (addra_pipe_1_net),
		.i0 (net_67),
		.i1 (net_78),
		.o (net_81)
	);
fifo2ram_emb_v1_AND u21 (
		.i0 (net_83),
		.i1 (net_82),
		.o (net_69)
	);
fifo2ram_emb_v1_AND u22 (
		.i0 (net_83),
		.i1 (ar[1]),
		.o (net_80)
	);
fifo2ram_emb_v1_NOT u23 (
		.i (ar[1]),
		.o (net_82)
	);
fifo2ram_emb_v1_ADDR_PIPE_A u_addra_pipe_2 (
		.clk (clkr),
		.ena (cer),
		.i (ar[2]),
		.o (addra_pipe_2_net)
	);
fifo2ram_emb_v1_MUX u24 (
		.sel (addra_pipe_2_net),
		.i0 (net_56),
		.i1 (net_81),
		.o (net_85)
	);
fifo2ram_emb_v1_AND u25 (
		.i0 (net_87),
		.i1 (net_86),
		.o (net_58)
	);
fifo2ram_emb_v1_AND u26 (
		.i0 (net_87),
		.i1 (ar[2]),
		.o (net_83)
	);
fifo2ram_emb_v1_NOT u27 (
		.i (ar[2]),
		.o (net_86)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_32 (
		.doa ({nc17137, nc17138, nc17139, nc17140, nc17141, nc17142, nc17143, nc17144, nc17145, nc17146, nc17147, nc17148, nc17149, nc17150, nc17151, nc17152, nc17153, nc17154, nc17155, nc17156, nc17157, nc17158, nc17159, nc17160, nc17161, nc17162, nc17163, nc17164, nc17165, nc17166, nc17167, nc17168, nc17169, nc17170, nc17171, nc17172, nc17173, nc17174, nc17175, nc17176, nc17177, nc17178, nc17179, nc17180, nc17181, nc17182, nc17183, nc17184, nc17185, nc17186, nc17187, nc17188, nc17189, nc17190, nc17191, nc17192, nc17193, nc17194, nc17195, nc17196, nc17197, nc17198, nc17199, net_90}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17200, nc17201, nc17202, nc17203, nc17204, nc17205, nc17206, nc17207, nc17208, nc17209, nc17210, nc17211, nc17212, nc17213, nc17214, nc17215, nc17216, nc17217, nc17218, nc17219, nc17220, nc17221, nc17222, nc17223, nc17224, nc17225, nc17226, nc17227, nc17228, nc17229, nc17230, nc17231, nc17232, nc17233, nc17234, nc17235, nc17236, nc17237, nc17238, nc17239, nc17240, nc17241, nc17242, nc17243, nc17244, nc17245, nc17246, nc17247, nc17248, nc17249, nc17250, nc17251, nc17252, nc17253, nc17254, nc17255, nc17256, nc17257, nc17258, nc17259, nc17260, nc17261, nc17262, dw[64]}),
		.dipa (),
		.dipb (),
		.cea (net_88),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_36 (
		.doa ({nc17263, nc17264, nc17265, nc17266, nc17267, nc17268, nc17269, nc17270, nc17271, nc17272, nc17273, nc17274, nc17275, nc17276, nc17277, nc17278, nc17279, nc17280, nc17281, nc17282, nc17283, nc17284, nc17285, nc17286, nc17287, nc17288, nc17289, nc17290, nc17291, nc17292, nc17293, nc17294, nc17295, nc17296, nc17297, nc17298, nc17299, nc17300, nc17301, nc17302, nc17303, nc17304, nc17305, nc17306, nc17307, nc17308, nc17309, nc17310, nc17311, nc17312, nc17313, nc17314, nc17315, nc17316, nc17317, nc17318, nc17319, nc17320, nc17321, nc17322, nc17323, nc17324, nc17325, net_94}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17326, nc17327, nc17328, nc17329, nc17330, nc17331, nc17332, nc17333, nc17334, nc17335, nc17336, nc17337, nc17338, nc17339, nc17340, nc17341, nc17342, nc17343, nc17344, nc17345, nc17346, nc17347, nc17348, nc17349, nc17350, nc17351, nc17352, nc17353, nc17354, nc17355, nc17356, nc17357, nc17358, nc17359, nc17360, nc17361, nc17362, nc17363, nc17364, nc17365, nc17366, nc17367, nc17368, nc17369, nc17370, nc17371, nc17372, nc17373, nc17374, nc17375, nc17376, nc17377, nc17378, nc17379, nc17380, nc17381, nc17382, nc17383, nc17384, nc17385, nc17386, nc17387, nc17388, dw[72]}),
		.dipa (),
		.dipb (),
		.cea (net_92),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u28 (
		.sel (addra_pipe_0_net),
		.i0 (net_90),
		.i1 (net_94),
		.o (net_96)
	);
fifo2ram_emb_v1_AND u29 (
		.i0 (net_98),
		.i1 (net_97),
		.o (net_88)
	);
fifo2ram_emb_v1_AND u30 (
		.i0 (net_98),
		.i1 (ar[0]),
		.o (net_92)
	);
fifo2ram_emb_v1_NOT u31 (
		.i (ar[0]),
		.o (net_97)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_40 (
		.doa ({nc17389, nc17390, nc17391, nc17392, nc17393, nc17394, nc17395, nc17396, nc17397, nc17398, nc17399, nc17400, nc17401, nc17402, nc17403, nc17404, nc17405, nc17406, nc17407, nc17408, nc17409, nc17410, nc17411, nc17412, nc17413, nc17414, nc17415, nc17416, nc17417, nc17418, nc17419, nc17420, nc17421, nc17422, nc17423, nc17424, nc17425, nc17426, nc17427, nc17428, nc17429, nc17430, nc17431, nc17432, nc17433, nc17434, nc17435, nc17436, nc17437, nc17438, nc17439, nc17440, nc17441, nc17442, nc17443, nc17444, nc17445, nc17446, nc17447, nc17448, nc17449, nc17450, nc17451, net_101}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17452, nc17453, nc17454, nc17455, nc17456, nc17457, nc17458, nc17459, nc17460, nc17461, nc17462, nc17463, nc17464, nc17465, nc17466, nc17467, nc17468, nc17469, nc17470, nc17471, nc17472, nc17473, nc17474, nc17475, nc17476, nc17477, nc17478, nc17479, nc17480, nc17481, nc17482, nc17483, nc17484, nc17485, nc17486, nc17487, nc17488, nc17489, nc17490, nc17491, nc17492, nc17493, nc17494, nc17495, nc17496, nc17497, nc17498, nc17499, nc17500, nc17501, nc17502, nc17503, nc17504, nc17505, nc17506, nc17507, nc17508, nc17509, nc17510, nc17511, nc17512, nc17513, nc17514, dw[80]}),
		.dipa (),
		.dipb (),
		.cea (net_99),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_44 (
		.doa ({nc17515, nc17516, nc17517, nc17518, nc17519, nc17520, nc17521, nc17522, nc17523, nc17524, nc17525, nc17526, nc17527, nc17528, nc17529, nc17530, nc17531, nc17532, nc17533, nc17534, nc17535, nc17536, nc17537, nc17538, nc17539, nc17540, nc17541, nc17542, nc17543, nc17544, nc17545, nc17546, nc17547, nc17548, nc17549, nc17550, nc17551, nc17552, nc17553, nc17554, nc17555, nc17556, nc17557, nc17558, nc17559, nc17560, nc17561, nc17562, nc17563, nc17564, nc17565, nc17566, nc17567, nc17568, nc17569, nc17570, nc17571, nc17572, nc17573, nc17574, nc17575, nc17576, nc17577, net_105}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17578, nc17579, nc17580, nc17581, nc17582, nc17583, nc17584, nc17585, nc17586, nc17587, nc17588, nc17589, nc17590, nc17591, nc17592, nc17593, nc17594, nc17595, nc17596, nc17597, nc17598, nc17599, nc17600, nc17601, nc17602, nc17603, nc17604, nc17605, nc17606, nc17607, nc17608, nc17609, nc17610, nc17611, nc17612, nc17613, nc17614, nc17615, nc17616, nc17617, nc17618, nc17619, nc17620, nc17621, nc17622, nc17623, nc17624, nc17625, nc17626, nc17627, nc17628, nc17629, nc17630, nc17631, nc17632, nc17633, nc17634, nc17635, nc17636, nc17637, nc17638, nc17639, nc17640, dw[88]}),
		.dipa (),
		.dipb (),
		.cea (net_103),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u32 (
		.sel (addra_pipe_0_net),
		.i0 (net_101),
		.i1 (net_105),
		.o (net_107)
	);
fifo2ram_emb_v1_AND u33 (
		.i0 (net_109),
		.i1 (net_108),
		.o (net_99)
	);
fifo2ram_emb_v1_AND u34 (
		.i0 (net_109),
		.i1 (ar[0]),
		.o (net_103)
	);
fifo2ram_emb_v1_NOT u35 (
		.i (ar[0]),
		.o (net_108)
	);
fifo2ram_emb_v1_MUX u36 (
		.sel (addra_pipe_1_net),
		.i0 (net_96),
		.i1 (net_107),
		.o (net_110)
	);
fifo2ram_emb_v1_AND u37 (
		.i0 (net_112),
		.i1 (net_111),
		.o (net_98)
	);
fifo2ram_emb_v1_AND u38 (
		.i0 (net_112),
		.i1 (ar[1]),
		.o (net_109)
	);
fifo2ram_emb_v1_NOT u39 (
		.i (ar[1]),
		.o (net_111)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_48 (
		.doa ({nc17641, nc17642, nc17643, nc17644, nc17645, nc17646, nc17647, nc17648, nc17649, nc17650, nc17651, nc17652, nc17653, nc17654, nc17655, nc17656, nc17657, nc17658, nc17659, nc17660, nc17661, nc17662, nc17663, nc17664, nc17665, nc17666, nc17667, nc17668, nc17669, nc17670, nc17671, nc17672, nc17673, nc17674, nc17675, nc17676, nc17677, nc17678, nc17679, nc17680, nc17681, nc17682, nc17683, nc17684, nc17685, nc17686, nc17687, nc17688, nc17689, nc17690, nc17691, nc17692, nc17693, nc17694, nc17695, nc17696, nc17697, nc17698, nc17699, nc17700, nc17701, nc17702, nc17703, net_115}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17704, nc17705, nc17706, nc17707, nc17708, nc17709, nc17710, nc17711, nc17712, nc17713, nc17714, nc17715, nc17716, nc17717, nc17718, nc17719, nc17720, nc17721, nc17722, nc17723, nc17724, nc17725, nc17726, nc17727, nc17728, nc17729, nc17730, nc17731, nc17732, nc17733, nc17734, nc17735, nc17736, nc17737, nc17738, nc17739, nc17740, nc17741, nc17742, nc17743, nc17744, nc17745, nc17746, nc17747, nc17748, nc17749, nc17750, nc17751, nc17752, nc17753, nc17754, nc17755, nc17756, nc17757, nc17758, nc17759, nc17760, nc17761, nc17762, nc17763, nc17764, nc17765, nc17766, dw[96]}),
		.dipa (),
		.dipb (),
		.cea (net_113),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_52 (
		.doa ({nc17767, nc17768, nc17769, nc17770, nc17771, nc17772, nc17773, nc17774, nc17775, nc17776, nc17777, nc17778, nc17779, nc17780, nc17781, nc17782, nc17783, nc17784, nc17785, nc17786, nc17787, nc17788, nc17789, nc17790, nc17791, nc17792, nc17793, nc17794, nc17795, nc17796, nc17797, nc17798, nc17799, nc17800, nc17801, nc17802, nc17803, nc17804, nc17805, nc17806, nc17807, nc17808, nc17809, nc17810, nc17811, nc17812, nc17813, nc17814, nc17815, nc17816, nc17817, nc17818, nc17819, nc17820, nc17821, nc17822, nc17823, nc17824, nc17825, nc17826, nc17827, nc17828, nc17829, net_119}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17830, nc17831, nc17832, nc17833, nc17834, nc17835, nc17836, nc17837, nc17838, nc17839, nc17840, nc17841, nc17842, nc17843, nc17844, nc17845, nc17846, nc17847, nc17848, nc17849, nc17850, nc17851, nc17852, nc17853, nc17854, nc17855, nc17856, nc17857, nc17858, nc17859, nc17860, nc17861, nc17862, nc17863, nc17864, nc17865, nc17866, nc17867, nc17868, nc17869, nc17870, nc17871, nc17872, nc17873, nc17874, nc17875, nc17876, nc17877, nc17878, nc17879, nc17880, nc17881, nc17882, nc17883, nc17884, nc17885, nc17886, nc17887, nc17888, nc17889, nc17890, nc17891, nc17892, dw[104]}),
		.dipa (),
		.dipb (),
		.cea (net_117),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u40 (
		.sel (addra_pipe_0_net),
		.i0 (net_115),
		.i1 (net_119),
		.o (net_121)
	);
fifo2ram_emb_v1_AND u41 (
		.i0 (net_123),
		.i1 (net_122),
		.o (net_113)
	);
fifo2ram_emb_v1_AND u42 (
		.i0 (net_123),
		.i1 (ar[0]),
		.o (net_117)
	);
fifo2ram_emb_v1_NOT u43 (
		.i (ar[0]),
		.o (net_122)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_56 (
		.doa ({nc17893, nc17894, nc17895, nc17896, nc17897, nc17898, nc17899, nc17900, nc17901, nc17902, nc17903, nc17904, nc17905, nc17906, nc17907, nc17908, nc17909, nc17910, nc17911, nc17912, nc17913, nc17914, nc17915, nc17916, nc17917, nc17918, nc17919, nc17920, nc17921, nc17922, nc17923, nc17924, nc17925, nc17926, nc17927, nc17928, nc17929, nc17930, nc17931, nc17932, nc17933, nc17934, nc17935, nc17936, nc17937, nc17938, nc17939, nc17940, nc17941, nc17942, nc17943, nc17944, nc17945, nc17946, nc17947, nc17948, nc17949, nc17950, nc17951, nc17952, nc17953, nc17954, nc17955, net_126}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc17956, nc17957, nc17958, nc17959, nc17960, nc17961, nc17962, nc17963, nc17964, nc17965, nc17966, nc17967, nc17968, nc17969, nc17970, nc17971, nc17972, nc17973, nc17974, nc17975, nc17976, nc17977, nc17978, nc17979, nc17980, nc17981, nc17982, nc17983, nc17984, nc17985, nc17986, nc17987, nc17988, nc17989, nc17990, nc17991, nc17992, nc17993, nc17994, nc17995, nc17996, nc17997, nc17998, nc17999, nc18000, nc18001, nc18002, nc18003, nc18004, nc18005, nc18006, nc18007, nc18008, nc18009, nc18010, nc18011, nc18012, nc18013, nc18014, nc18015, nc18016, nc18017, nc18018, dw[112]}),
		.dipa (),
		.dipb (),
		.cea (net_124),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_60 (
		.doa ({nc18019, nc18020, nc18021, nc18022, nc18023, nc18024, nc18025, nc18026, nc18027, nc18028, nc18029, nc18030, nc18031, nc18032, nc18033, nc18034, nc18035, nc18036, nc18037, nc18038, nc18039, nc18040, nc18041, nc18042, nc18043, nc18044, nc18045, nc18046, nc18047, nc18048, nc18049, nc18050, nc18051, nc18052, nc18053, nc18054, nc18055, nc18056, nc18057, nc18058, nc18059, nc18060, nc18061, nc18062, nc18063, nc18064, nc18065, nc18066, nc18067, nc18068, nc18069, nc18070, nc18071, nc18072, nc18073, nc18074, nc18075, nc18076, nc18077, nc18078, nc18079, nc18080, nc18081, net_130}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18082, nc18083, nc18084, nc18085, nc18086, nc18087, nc18088, nc18089, nc18090, nc18091, nc18092, nc18093, nc18094, nc18095, nc18096, nc18097, nc18098, nc18099, nc18100, nc18101, nc18102, nc18103, nc18104, nc18105, nc18106, nc18107, nc18108, nc18109, nc18110, nc18111, nc18112, nc18113, nc18114, nc18115, nc18116, nc18117, nc18118, nc18119, nc18120, nc18121, nc18122, nc18123, nc18124, nc18125, nc18126, nc18127, nc18128, nc18129, nc18130, nc18131, nc18132, nc18133, nc18134, nc18135, nc18136, nc18137, nc18138, nc18139, nc18140, nc18141, nc18142, nc18143, nc18144, dw[120]}),
		.dipa (),
		.dipb (),
		.cea (net_128),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u44 (
		.sel (addra_pipe_0_net),
		.i0 (net_126),
		.i1 (net_130),
		.o (net_132)
	);
fifo2ram_emb_v1_AND u45 (
		.i0 (net_134),
		.i1 (net_133),
		.o (net_124)
	);
fifo2ram_emb_v1_AND u46 (
		.i0 (net_134),
		.i1 (ar[0]),
		.o (net_128)
	);
fifo2ram_emb_v1_NOT u47 (
		.i (ar[0]),
		.o (net_133)
	);
fifo2ram_emb_v1_MUX u48 (
		.sel (addra_pipe_1_net),
		.i0 (net_121),
		.i1 (net_132),
		.o (net_135)
	);
fifo2ram_emb_v1_AND u49 (
		.i0 (net_137),
		.i1 (net_136),
		.o (net_123)
	);
fifo2ram_emb_v1_AND u50 (
		.i0 (net_137),
		.i1 (ar[1]),
		.o (net_134)
	);
fifo2ram_emb_v1_NOT u51 (
		.i (ar[1]),
		.o (net_136)
	);
fifo2ram_emb_v1_MUX u52 (
		.sel (addra_pipe_2_net),
		.i0 (net_110),
		.i1 (net_135),
		.o (net_138)
	);
fifo2ram_emb_v1_AND u53 (
		.i0 (net_140),
		.i1 (net_139),
		.o (net_112)
	);
fifo2ram_emb_v1_AND u54 (
		.i0 (net_140),
		.i1 (ar[2]),
		.o (net_137)
	);
fifo2ram_emb_v1_NOT u55 (
		.i (ar[2]),
		.o (net_139)
	);
fifo2ram_emb_v1_ADDR_PIPE_A u_addra_pipe_3 (
		.clk (clkr),
		.ena (cer),
		.i (ar[3]),
		.o (addra_pipe_3_net)
	);
fifo2ram_emb_v1_MUX u56 (
		.sel (addra_pipe_3_net),
		.i0 (net_85),
		.i1 (net_138),
		.o (qr[0])
	);
fifo2ram_emb_v1_AND u57 (
		.i0 (cer),
		.i1 (net_143),
		.o (net_87)
	);
fifo2ram_emb_v1_AND u58 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_140)
	);
fifo2ram_emb_v1_NOT u59 (
		.i (ar[3]),
		.o (net_143)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_64 (
		.doa ({nc18145, nc18146, nc18147, nc18148, nc18149, nc18150, nc18151, nc18152, nc18153, nc18154, nc18155, nc18156, nc18157, nc18158, nc18159, nc18160, nc18161, nc18162, nc18163, nc18164, nc18165, nc18166, nc18167, nc18168, nc18169, nc18170, nc18171, nc18172, nc18173, nc18174, nc18175, nc18176, nc18177, nc18178, nc18179, nc18180, nc18181, nc18182, nc18183, nc18184, nc18185, nc18186, nc18187, nc18188, nc18189, nc18190, nc18191, nc18192, nc18193, nc18194, nc18195, nc18196, nc18197, nc18198, nc18199, nc18200, nc18201, nc18202, nc18203, nc18204, nc18205, nc18206, nc18207, net_147}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18208, nc18209, nc18210, nc18211, nc18212, nc18213, nc18214, nc18215, nc18216, nc18217, nc18218, nc18219, nc18220, nc18221, nc18222, nc18223, nc18224, nc18225, nc18226, nc18227, nc18228, nc18229, nc18230, nc18231, nc18232, nc18233, nc18234, nc18235, nc18236, nc18237, nc18238, nc18239, nc18240, nc18241, nc18242, nc18243, nc18244, nc18245, nc18246, nc18247, nc18248, nc18249, nc18250, nc18251, nc18252, nc18253, nc18254, nc18255, nc18256, nc18257, nc18258, nc18259, nc18260, nc18261, nc18262, nc18263, nc18264, nc18265, nc18266, nc18267, nc18268, nc18269, nc18270, dw[1]}),
		.dipa (),
		.dipb (),
		.cea (net_145),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_68 (
		.doa ({nc18271, nc18272, nc18273, nc18274, nc18275, nc18276, nc18277, nc18278, nc18279, nc18280, nc18281, nc18282, nc18283, nc18284, nc18285, nc18286, nc18287, nc18288, nc18289, nc18290, nc18291, nc18292, nc18293, nc18294, nc18295, nc18296, nc18297, nc18298, nc18299, nc18300, nc18301, nc18302, nc18303, nc18304, nc18305, nc18306, nc18307, nc18308, nc18309, nc18310, nc18311, nc18312, nc18313, nc18314, nc18315, nc18316, nc18317, nc18318, nc18319, nc18320, nc18321, nc18322, nc18323, nc18324, nc18325, nc18326, nc18327, nc18328, nc18329, nc18330, nc18331, nc18332, nc18333, net_151}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18334, nc18335, nc18336, nc18337, nc18338, nc18339, nc18340, nc18341, nc18342, nc18343, nc18344, nc18345, nc18346, nc18347, nc18348, nc18349, nc18350, nc18351, nc18352, nc18353, nc18354, nc18355, nc18356, nc18357, nc18358, nc18359, nc18360, nc18361, nc18362, nc18363, nc18364, nc18365, nc18366, nc18367, nc18368, nc18369, nc18370, nc18371, nc18372, nc18373, nc18374, nc18375, nc18376, nc18377, nc18378, nc18379, nc18380, nc18381, nc18382, nc18383, nc18384, nc18385, nc18386, nc18387, nc18388, nc18389, nc18390, nc18391, nc18392, nc18393, nc18394, nc18395, nc18396, dw[9]}),
		.dipa (),
		.dipb (),
		.cea (net_149),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u60 (
		.sel (addra_pipe_0_net),
		.i0 (net_147),
		.i1 (net_151),
		.o (net_153)
	);
fifo2ram_emb_v1_AND u61 (
		.i0 (net_155),
		.i1 (net_154),
		.o (net_145)
	);
fifo2ram_emb_v1_AND u62 (
		.i0 (net_155),
		.i1 (ar[0]),
		.o (net_149)
	);
fifo2ram_emb_v1_NOT u63 (
		.i (ar[0]),
		.o (net_154)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_72 (
		.doa ({nc18397, nc18398, nc18399, nc18400, nc18401, nc18402, nc18403, nc18404, nc18405, nc18406, nc18407, nc18408, nc18409, nc18410, nc18411, nc18412, nc18413, nc18414, nc18415, nc18416, nc18417, nc18418, nc18419, nc18420, nc18421, nc18422, nc18423, nc18424, nc18425, nc18426, nc18427, nc18428, nc18429, nc18430, nc18431, nc18432, nc18433, nc18434, nc18435, nc18436, nc18437, nc18438, nc18439, nc18440, nc18441, nc18442, nc18443, nc18444, nc18445, nc18446, nc18447, nc18448, nc18449, nc18450, nc18451, nc18452, nc18453, nc18454, nc18455, nc18456, nc18457, nc18458, nc18459, net_158}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18460, nc18461, nc18462, nc18463, nc18464, nc18465, nc18466, nc18467, nc18468, nc18469, nc18470, nc18471, nc18472, nc18473, nc18474, nc18475, nc18476, nc18477, nc18478, nc18479, nc18480, nc18481, nc18482, nc18483, nc18484, nc18485, nc18486, nc18487, nc18488, nc18489, nc18490, nc18491, nc18492, nc18493, nc18494, nc18495, nc18496, nc18497, nc18498, nc18499, nc18500, nc18501, nc18502, nc18503, nc18504, nc18505, nc18506, nc18507, nc18508, nc18509, nc18510, nc18511, nc18512, nc18513, nc18514, nc18515, nc18516, nc18517, nc18518, nc18519, nc18520, nc18521, nc18522, dw[17]}),
		.dipa (),
		.dipb (),
		.cea (net_156),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_76 (
		.doa ({nc18523, nc18524, nc18525, nc18526, nc18527, nc18528, nc18529, nc18530, nc18531, nc18532, nc18533, nc18534, nc18535, nc18536, nc18537, nc18538, nc18539, nc18540, nc18541, nc18542, nc18543, nc18544, nc18545, nc18546, nc18547, nc18548, nc18549, nc18550, nc18551, nc18552, nc18553, nc18554, nc18555, nc18556, nc18557, nc18558, nc18559, nc18560, nc18561, nc18562, nc18563, nc18564, nc18565, nc18566, nc18567, nc18568, nc18569, nc18570, nc18571, nc18572, nc18573, nc18574, nc18575, nc18576, nc18577, nc18578, nc18579, nc18580, nc18581, nc18582, nc18583, nc18584, nc18585, net_162}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18586, nc18587, nc18588, nc18589, nc18590, nc18591, nc18592, nc18593, nc18594, nc18595, nc18596, nc18597, nc18598, nc18599, nc18600, nc18601, nc18602, nc18603, nc18604, nc18605, nc18606, nc18607, nc18608, nc18609, nc18610, nc18611, nc18612, nc18613, nc18614, nc18615, nc18616, nc18617, nc18618, nc18619, nc18620, nc18621, nc18622, nc18623, nc18624, nc18625, nc18626, nc18627, nc18628, nc18629, nc18630, nc18631, nc18632, nc18633, nc18634, nc18635, nc18636, nc18637, nc18638, nc18639, nc18640, nc18641, nc18642, nc18643, nc18644, nc18645, nc18646, nc18647, nc18648, dw[25]}),
		.dipa (),
		.dipb (),
		.cea (net_160),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u64 (
		.sel (addra_pipe_0_net),
		.i0 (net_158),
		.i1 (net_162),
		.o (net_164)
	);
fifo2ram_emb_v1_AND u65 (
		.i0 (net_166),
		.i1 (net_165),
		.o (net_156)
	);
fifo2ram_emb_v1_AND u66 (
		.i0 (net_166),
		.i1 (ar[0]),
		.o (net_160)
	);
fifo2ram_emb_v1_NOT u67 (
		.i (ar[0]),
		.o (net_165)
	);
fifo2ram_emb_v1_MUX u68 (
		.sel (addra_pipe_1_net),
		.i0 (net_153),
		.i1 (net_164),
		.o (net_167)
	);
fifo2ram_emb_v1_AND u69 (
		.i0 (net_169),
		.i1 (net_168),
		.o (net_155)
	);
fifo2ram_emb_v1_AND u70 (
		.i0 (net_169),
		.i1 (ar[1]),
		.o (net_166)
	);
fifo2ram_emb_v1_NOT u71 (
		.i (ar[1]),
		.o (net_168)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_80 (
		.doa ({nc18649, nc18650, nc18651, nc18652, nc18653, nc18654, nc18655, nc18656, nc18657, nc18658, nc18659, nc18660, nc18661, nc18662, nc18663, nc18664, nc18665, nc18666, nc18667, nc18668, nc18669, nc18670, nc18671, nc18672, nc18673, nc18674, nc18675, nc18676, nc18677, nc18678, nc18679, nc18680, nc18681, nc18682, nc18683, nc18684, nc18685, nc18686, nc18687, nc18688, nc18689, nc18690, nc18691, nc18692, nc18693, nc18694, nc18695, nc18696, nc18697, nc18698, nc18699, nc18700, nc18701, nc18702, nc18703, nc18704, nc18705, nc18706, nc18707, nc18708, nc18709, nc18710, nc18711, net_172}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18712, nc18713, nc18714, nc18715, nc18716, nc18717, nc18718, nc18719, nc18720, nc18721, nc18722, nc18723, nc18724, nc18725, nc18726, nc18727, nc18728, nc18729, nc18730, nc18731, nc18732, nc18733, nc18734, nc18735, nc18736, nc18737, nc18738, nc18739, nc18740, nc18741, nc18742, nc18743, nc18744, nc18745, nc18746, nc18747, nc18748, nc18749, nc18750, nc18751, nc18752, nc18753, nc18754, nc18755, nc18756, nc18757, nc18758, nc18759, nc18760, nc18761, nc18762, nc18763, nc18764, nc18765, nc18766, nc18767, nc18768, nc18769, nc18770, nc18771, nc18772, nc18773, nc18774, dw[33]}),
		.dipa (),
		.dipb (),
		.cea (net_170),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_84 (
		.doa ({nc18775, nc18776, nc18777, nc18778, nc18779, nc18780, nc18781, nc18782, nc18783, nc18784, nc18785, nc18786, nc18787, nc18788, nc18789, nc18790, nc18791, nc18792, nc18793, nc18794, nc18795, nc18796, nc18797, nc18798, nc18799, nc18800, nc18801, nc18802, nc18803, nc18804, nc18805, nc18806, nc18807, nc18808, nc18809, nc18810, nc18811, nc18812, nc18813, nc18814, nc18815, nc18816, nc18817, nc18818, nc18819, nc18820, nc18821, nc18822, nc18823, nc18824, nc18825, nc18826, nc18827, nc18828, nc18829, nc18830, nc18831, nc18832, nc18833, nc18834, nc18835, nc18836, nc18837, net_176}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18838, nc18839, nc18840, nc18841, nc18842, nc18843, nc18844, nc18845, nc18846, nc18847, nc18848, nc18849, nc18850, nc18851, nc18852, nc18853, nc18854, nc18855, nc18856, nc18857, nc18858, nc18859, nc18860, nc18861, nc18862, nc18863, nc18864, nc18865, nc18866, nc18867, nc18868, nc18869, nc18870, nc18871, nc18872, nc18873, nc18874, nc18875, nc18876, nc18877, nc18878, nc18879, nc18880, nc18881, nc18882, nc18883, nc18884, nc18885, nc18886, nc18887, nc18888, nc18889, nc18890, nc18891, nc18892, nc18893, nc18894, nc18895, nc18896, nc18897, nc18898, nc18899, nc18900, dw[41]}),
		.dipa (),
		.dipb (),
		.cea (net_174),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u72 (
		.sel (addra_pipe_0_net),
		.i0 (net_172),
		.i1 (net_176),
		.o (net_178)
	);
fifo2ram_emb_v1_AND u73 (
		.i0 (net_180),
		.i1 (net_179),
		.o (net_170)
	);
fifo2ram_emb_v1_AND u74 (
		.i0 (net_180),
		.i1 (ar[0]),
		.o (net_174)
	);
fifo2ram_emb_v1_NOT u75 (
		.i (ar[0]),
		.o (net_179)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_88 (
		.doa ({nc18901, nc18902, nc18903, nc18904, nc18905, nc18906, nc18907, nc18908, nc18909, nc18910, nc18911, nc18912, nc18913, nc18914, nc18915, nc18916, nc18917, nc18918, nc18919, nc18920, nc18921, nc18922, nc18923, nc18924, nc18925, nc18926, nc18927, nc18928, nc18929, nc18930, nc18931, nc18932, nc18933, nc18934, nc18935, nc18936, nc18937, nc18938, nc18939, nc18940, nc18941, nc18942, nc18943, nc18944, nc18945, nc18946, nc18947, nc18948, nc18949, nc18950, nc18951, nc18952, nc18953, nc18954, nc18955, nc18956, nc18957, nc18958, nc18959, nc18960, nc18961, nc18962, nc18963, net_183}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc18964, nc18965, nc18966, nc18967, nc18968, nc18969, nc18970, nc18971, nc18972, nc18973, nc18974, nc18975, nc18976, nc18977, nc18978, nc18979, nc18980, nc18981, nc18982, nc18983, nc18984, nc18985, nc18986, nc18987, nc18988, nc18989, nc18990, nc18991, nc18992, nc18993, nc18994, nc18995, nc18996, nc18997, nc18998, nc18999, nc19000, nc19001, nc19002, nc19003, nc19004, nc19005, nc19006, nc19007, nc19008, nc19009, nc19010, nc19011, nc19012, nc19013, nc19014, nc19015, nc19016, nc19017, nc19018, nc19019, nc19020, nc19021, nc19022, nc19023, nc19024, nc19025, nc19026, dw[49]}),
		.dipa (),
		.dipb (),
		.cea (net_181),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_92 (
		.doa ({nc19027, nc19028, nc19029, nc19030, nc19031, nc19032, nc19033, nc19034, nc19035, nc19036, nc19037, nc19038, nc19039, nc19040, nc19041, nc19042, nc19043, nc19044, nc19045, nc19046, nc19047, nc19048, nc19049, nc19050, nc19051, nc19052, nc19053, nc19054, nc19055, nc19056, nc19057, nc19058, nc19059, nc19060, nc19061, nc19062, nc19063, nc19064, nc19065, nc19066, nc19067, nc19068, nc19069, nc19070, nc19071, nc19072, nc19073, nc19074, nc19075, nc19076, nc19077, nc19078, nc19079, nc19080, nc19081, nc19082, nc19083, nc19084, nc19085, nc19086, nc19087, nc19088, nc19089, net_187}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19090, nc19091, nc19092, nc19093, nc19094, nc19095, nc19096, nc19097, nc19098, nc19099, nc19100, nc19101, nc19102, nc19103, nc19104, nc19105, nc19106, nc19107, nc19108, nc19109, nc19110, nc19111, nc19112, nc19113, nc19114, nc19115, nc19116, nc19117, nc19118, nc19119, nc19120, nc19121, nc19122, nc19123, nc19124, nc19125, nc19126, nc19127, nc19128, nc19129, nc19130, nc19131, nc19132, nc19133, nc19134, nc19135, nc19136, nc19137, nc19138, nc19139, nc19140, nc19141, nc19142, nc19143, nc19144, nc19145, nc19146, nc19147, nc19148, nc19149, nc19150, nc19151, nc19152, dw[57]}),
		.dipa (),
		.dipb (),
		.cea (net_185),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u76 (
		.sel (addra_pipe_0_net),
		.i0 (net_183),
		.i1 (net_187),
		.o (net_189)
	);
fifo2ram_emb_v1_AND u77 (
		.i0 (net_191),
		.i1 (net_190),
		.o (net_181)
	);
fifo2ram_emb_v1_AND u78 (
		.i0 (net_191),
		.i1 (ar[0]),
		.o (net_185)
	);
fifo2ram_emb_v1_NOT u79 (
		.i (ar[0]),
		.o (net_190)
	);
fifo2ram_emb_v1_MUX u80 (
		.sel (addra_pipe_1_net),
		.i0 (net_178),
		.i1 (net_189),
		.o (net_192)
	);
fifo2ram_emb_v1_AND u81 (
		.i0 (net_194),
		.i1 (net_193),
		.o (net_180)
	);
fifo2ram_emb_v1_AND u82 (
		.i0 (net_194),
		.i1 (ar[1]),
		.o (net_191)
	);
fifo2ram_emb_v1_NOT u83 (
		.i (ar[1]),
		.o (net_193)
	);
fifo2ram_emb_v1_MUX u84 (
		.sel (addra_pipe_2_net),
		.i0 (net_167),
		.i1 (net_192),
		.o (net_195)
	);
fifo2ram_emb_v1_AND u85 (
		.i0 (net_197),
		.i1 (net_196),
		.o (net_169)
	);
fifo2ram_emb_v1_AND u86 (
		.i0 (net_197),
		.i1 (ar[2]),
		.o (net_194)
	);
fifo2ram_emb_v1_NOT u87 (
		.i (ar[2]),
		.o (net_196)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_96 (
		.doa ({nc19153, nc19154, nc19155, nc19156, nc19157, nc19158, nc19159, nc19160, nc19161, nc19162, nc19163, nc19164, nc19165, nc19166, nc19167, nc19168, nc19169, nc19170, nc19171, nc19172, nc19173, nc19174, nc19175, nc19176, nc19177, nc19178, nc19179, nc19180, nc19181, nc19182, nc19183, nc19184, nc19185, nc19186, nc19187, nc19188, nc19189, nc19190, nc19191, nc19192, nc19193, nc19194, nc19195, nc19196, nc19197, nc19198, nc19199, nc19200, nc19201, nc19202, nc19203, nc19204, nc19205, nc19206, nc19207, nc19208, nc19209, nc19210, nc19211, nc19212, nc19213, nc19214, nc19215, net_200}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19216, nc19217, nc19218, nc19219, nc19220, nc19221, nc19222, nc19223, nc19224, nc19225, nc19226, nc19227, nc19228, nc19229, nc19230, nc19231, nc19232, nc19233, nc19234, nc19235, nc19236, nc19237, nc19238, nc19239, nc19240, nc19241, nc19242, nc19243, nc19244, nc19245, nc19246, nc19247, nc19248, nc19249, nc19250, nc19251, nc19252, nc19253, nc19254, nc19255, nc19256, nc19257, nc19258, nc19259, nc19260, nc19261, nc19262, nc19263, nc19264, nc19265, nc19266, nc19267, nc19268, nc19269, nc19270, nc19271, nc19272, nc19273, nc19274, nc19275, nc19276, nc19277, nc19278, dw[65]}),
		.dipa (),
		.dipb (),
		.cea (net_198),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_100 (
		.doa ({nc19279, nc19280, nc19281, nc19282, nc19283, nc19284, nc19285, nc19286, nc19287, nc19288, nc19289, nc19290, nc19291, nc19292, nc19293, nc19294, nc19295, nc19296, nc19297, nc19298, nc19299, nc19300, nc19301, nc19302, nc19303, nc19304, nc19305, nc19306, nc19307, nc19308, nc19309, nc19310, nc19311, nc19312, nc19313, nc19314, nc19315, nc19316, nc19317, nc19318, nc19319, nc19320, nc19321, nc19322, nc19323, nc19324, nc19325, nc19326, nc19327, nc19328, nc19329, nc19330, nc19331, nc19332, nc19333, nc19334, nc19335, nc19336, nc19337, nc19338, nc19339, nc19340, nc19341, net_204}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19342, nc19343, nc19344, nc19345, nc19346, nc19347, nc19348, nc19349, nc19350, nc19351, nc19352, nc19353, nc19354, nc19355, nc19356, nc19357, nc19358, nc19359, nc19360, nc19361, nc19362, nc19363, nc19364, nc19365, nc19366, nc19367, nc19368, nc19369, nc19370, nc19371, nc19372, nc19373, nc19374, nc19375, nc19376, nc19377, nc19378, nc19379, nc19380, nc19381, nc19382, nc19383, nc19384, nc19385, nc19386, nc19387, nc19388, nc19389, nc19390, nc19391, nc19392, nc19393, nc19394, nc19395, nc19396, nc19397, nc19398, nc19399, nc19400, nc19401, nc19402, nc19403, nc19404, dw[73]}),
		.dipa (),
		.dipb (),
		.cea (net_202),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u88 (
		.sel (addra_pipe_0_net),
		.i0 (net_200),
		.i1 (net_204),
		.o (net_206)
	);
fifo2ram_emb_v1_AND u89 (
		.i0 (net_208),
		.i1 (net_207),
		.o (net_198)
	);
fifo2ram_emb_v1_AND u90 (
		.i0 (net_208),
		.i1 (ar[0]),
		.o (net_202)
	);
fifo2ram_emb_v1_NOT u91 (
		.i (ar[0]),
		.o (net_207)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_104 (
		.doa ({nc19405, nc19406, nc19407, nc19408, nc19409, nc19410, nc19411, nc19412, nc19413, nc19414, nc19415, nc19416, nc19417, nc19418, nc19419, nc19420, nc19421, nc19422, nc19423, nc19424, nc19425, nc19426, nc19427, nc19428, nc19429, nc19430, nc19431, nc19432, nc19433, nc19434, nc19435, nc19436, nc19437, nc19438, nc19439, nc19440, nc19441, nc19442, nc19443, nc19444, nc19445, nc19446, nc19447, nc19448, nc19449, nc19450, nc19451, nc19452, nc19453, nc19454, nc19455, nc19456, nc19457, nc19458, nc19459, nc19460, nc19461, nc19462, nc19463, nc19464, nc19465, nc19466, nc19467, net_211}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19468, nc19469, nc19470, nc19471, nc19472, nc19473, nc19474, nc19475, nc19476, nc19477, nc19478, nc19479, nc19480, nc19481, nc19482, nc19483, nc19484, nc19485, nc19486, nc19487, nc19488, nc19489, nc19490, nc19491, nc19492, nc19493, nc19494, nc19495, nc19496, nc19497, nc19498, nc19499, nc19500, nc19501, nc19502, nc19503, nc19504, nc19505, nc19506, nc19507, nc19508, nc19509, nc19510, nc19511, nc19512, nc19513, nc19514, nc19515, nc19516, nc19517, nc19518, nc19519, nc19520, nc19521, nc19522, nc19523, nc19524, nc19525, nc19526, nc19527, nc19528, nc19529, nc19530, dw[81]}),
		.dipa (),
		.dipb (),
		.cea (net_209),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_108 (
		.doa ({nc19531, nc19532, nc19533, nc19534, nc19535, nc19536, nc19537, nc19538, nc19539, nc19540, nc19541, nc19542, nc19543, nc19544, nc19545, nc19546, nc19547, nc19548, nc19549, nc19550, nc19551, nc19552, nc19553, nc19554, nc19555, nc19556, nc19557, nc19558, nc19559, nc19560, nc19561, nc19562, nc19563, nc19564, nc19565, nc19566, nc19567, nc19568, nc19569, nc19570, nc19571, nc19572, nc19573, nc19574, nc19575, nc19576, nc19577, nc19578, nc19579, nc19580, nc19581, nc19582, nc19583, nc19584, nc19585, nc19586, nc19587, nc19588, nc19589, nc19590, nc19591, nc19592, nc19593, net_215}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19594, nc19595, nc19596, nc19597, nc19598, nc19599, nc19600, nc19601, nc19602, nc19603, nc19604, nc19605, nc19606, nc19607, nc19608, nc19609, nc19610, nc19611, nc19612, nc19613, nc19614, nc19615, nc19616, nc19617, nc19618, nc19619, nc19620, nc19621, nc19622, nc19623, nc19624, nc19625, nc19626, nc19627, nc19628, nc19629, nc19630, nc19631, nc19632, nc19633, nc19634, nc19635, nc19636, nc19637, nc19638, nc19639, nc19640, nc19641, nc19642, nc19643, nc19644, nc19645, nc19646, nc19647, nc19648, nc19649, nc19650, nc19651, nc19652, nc19653, nc19654, nc19655, nc19656, dw[89]}),
		.dipa (),
		.dipb (),
		.cea (net_213),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u92 (
		.sel (addra_pipe_0_net),
		.i0 (net_211),
		.i1 (net_215),
		.o (net_217)
	);
fifo2ram_emb_v1_AND u93 (
		.i0 (net_219),
		.i1 (net_218),
		.o (net_209)
	);
fifo2ram_emb_v1_AND u94 (
		.i0 (net_219),
		.i1 (ar[0]),
		.o (net_213)
	);
fifo2ram_emb_v1_NOT u95 (
		.i (ar[0]),
		.o (net_218)
	);
fifo2ram_emb_v1_MUX u96 (
		.sel (addra_pipe_1_net),
		.i0 (net_206),
		.i1 (net_217),
		.o (net_220)
	);
fifo2ram_emb_v1_AND u97 (
		.i0 (net_222),
		.i1 (net_221),
		.o (net_208)
	);
fifo2ram_emb_v1_AND u98 (
		.i0 (net_222),
		.i1 (ar[1]),
		.o (net_219)
	);
fifo2ram_emb_v1_NOT u99 (
		.i (ar[1]),
		.o (net_221)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_112 (
		.doa ({nc19657, nc19658, nc19659, nc19660, nc19661, nc19662, nc19663, nc19664, nc19665, nc19666, nc19667, nc19668, nc19669, nc19670, nc19671, nc19672, nc19673, nc19674, nc19675, nc19676, nc19677, nc19678, nc19679, nc19680, nc19681, nc19682, nc19683, nc19684, nc19685, nc19686, nc19687, nc19688, nc19689, nc19690, nc19691, nc19692, nc19693, nc19694, nc19695, nc19696, nc19697, nc19698, nc19699, nc19700, nc19701, nc19702, nc19703, nc19704, nc19705, nc19706, nc19707, nc19708, nc19709, nc19710, nc19711, nc19712, nc19713, nc19714, nc19715, nc19716, nc19717, nc19718, nc19719, net_225}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19720, nc19721, nc19722, nc19723, nc19724, nc19725, nc19726, nc19727, nc19728, nc19729, nc19730, nc19731, nc19732, nc19733, nc19734, nc19735, nc19736, nc19737, nc19738, nc19739, nc19740, nc19741, nc19742, nc19743, nc19744, nc19745, nc19746, nc19747, nc19748, nc19749, nc19750, nc19751, nc19752, nc19753, nc19754, nc19755, nc19756, nc19757, nc19758, nc19759, nc19760, nc19761, nc19762, nc19763, nc19764, nc19765, nc19766, nc19767, nc19768, nc19769, nc19770, nc19771, nc19772, nc19773, nc19774, nc19775, nc19776, nc19777, nc19778, nc19779, nc19780, nc19781, nc19782, dw[97]}),
		.dipa (),
		.dipb (),
		.cea (net_223),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_116 (
		.doa ({nc19783, nc19784, nc19785, nc19786, nc19787, nc19788, nc19789, nc19790, nc19791, nc19792, nc19793, nc19794, nc19795, nc19796, nc19797, nc19798, nc19799, nc19800, nc19801, nc19802, nc19803, nc19804, nc19805, nc19806, nc19807, nc19808, nc19809, nc19810, nc19811, nc19812, nc19813, nc19814, nc19815, nc19816, nc19817, nc19818, nc19819, nc19820, nc19821, nc19822, nc19823, nc19824, nc19825, nc19826, nc19827, nc19828, nc19829, nc19830, nc19831, nc19832, nc19833, nc19834, nc19835, nc19836, nc19837, nc19838, nc19839, nc19840, nc19841, nc19842, nc19843, nc19844, nc19845, net_229}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19846, nc19847, nc19848, nc19849, nc19850, nc19851, nc19852, nc19853, nc19854, nc19855, nc19856, nc19857, nc19858, nc19859, nc19860, nc19861, nc19862, nc19863, nc19864, nc19865, nc19866, nc19867, nc19868, nc19869, nc19870, nc19871, nc19872, nc19873, nc19874, nc19875, nc19876, nc19877, nc19878, nc19879, nc19880, nc19881, nc19882, nc19883, nc19884, nc19885, nc19886, nc19887, nc19888, nc19889, nc19890, nc19891, nc19892, nc19893, nc19894, nc19895, nc19896, nc19897, nc19898, nc19899, nc19900, nc19901, nc19902, nc19903, nc19904, nc19905, nc19906, nc19907, nc19908, dw[105]}),
		.dipa (),
		.dipb (),
		.cea (net_227),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u100 (
		.sel (addra_pipe_0_net),
		.i0 (net_225),
		.i1 (net_229),
		.o (net_231)
	);
fifo2ram_emb_v1_AND u101 (
		.i0 (net_233),
		.i1 (net_232),
		.o (net_223)
	);
fifo2ram_emb_v1_AND u102 (
		.i0 (net_233),
		.i1 (ar[0]),
		.o (net_227)
	);
fifo2ram_emb_v1_NOT u103 (
		.i (ar[0]),
		.o (net_232)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_120 (
		.doa ({nc19909, nc19910, nc19911, nc19912, nc19913, nc19914, nc19915, nc19916, nc19917, nc19918, nc19919, nc19920, nc19921, nc19922, nc19923, nc19924, nc19925, nc19926, nc19927, nc19928, nc19929, nc19930, nc19931, nc19932, nc19933, nc19934, nc19935, nc19936, nc19937, nc19938, nc19939, nc19940, nc19941, nc19942, nc19943, nc19944, nc19945, nc19946, nc19947, nc19948, nc19949, nc19950, nc19951, nc19952, nc19953, nc19954, nc19955, nc19956, nc19957, nc19958, nc19959, nc19960, nc19961, nc19962, nc19963, nc19964, nc19965, nc19966, nc19967, nc19968, nc19969, nc19970, nc19971, net_236}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc19972, nc19973, nc19974, nc19975, nc19976, nc19977, nc19978, nc19979, nc19980, nc19981, nc19982, nc19983, nc19984, nc19985, nc19986, nc19987, nc19988, nc19989, nc19990, nc19991, nc19992, nc19993, nc19994, nc19995, nc19996, nc19997, nc19998, nc19999, nc20000, nc20001, nc20002, nc20003, nc20004, nc20005, nc20006, nc20007, nc20008, nc20009, nc20010, nc20011, nc20012, nc20013, nc20014, nc20015, nc20016, nc20017, nc20018, nc20019, nc20020, nc20021, nc20022, nc20023, nc20024, nc20025, nc20026, nc20027, nc20028, nc20029, nc20030, nc20031, nc20032, nc20033, nc20034, dw[113]}),
		.dipa (),
		.dipb (),
		.cea (net_234),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_124 (
		.doa ({nc20035, nc20036, nc20037, nc20038, nc20039, nc20040, nc20041, nc20042, nc20043, nc20044, nc20045, nc20046, nc20047, nc20048, nc20049, nc20050, nc20051, nc20052, nc20053, nc20054, nc20055, nc20056, nc20057, nc20058, nc20059, nc20060, nc20061, nc20062, nc20063, nc20064, nc20065, nc20066, nc20067, nc20068, nc20069, nc20070, nc20071, nc20072, nc20073, nc20074, nc20075, nc20076, nc20077, nc20078, nc20079, nc20080, nc20081, nc20082, nc20083, nc20084, nc20085, nc20086, nc20087, nc20088, nc20089, nc20090, nc20091, nc20092, nc20093, nc20094, nc20095, nc20096, nc20097, net_240}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20098, nc20099, nc20100, nc20101, nc20102, nc20103, nc20104, nc20105, nc20106, nc20107, nc20108, nc20109, nc20110, nc20111, nc20112, nc20113, nc20114, nc20115, nc20116, nc20117, nc20118, nc20119, nc20120, nc20121, nc20122, nc20123, nc20124, nc20125, nc20126, nc20127, nc20128, nc20129, nc20130, nc20131, nc20132, nc20133, nc20134, nc20135, nc20136, nc20137, nc20138, nc20139, nc20140, nc20141, nc20142, nc20143, nc20144, nc20145, nc20146, nc20147, nc20148, nc20149, nc20150, nc20151, nc20152, nc20153, nc20154, nc20155, nc20156, nc20157, nc20158, nc20159, nc20160, dw[121]}),
		.dipa (),
		.dipb (),
		.cea (net_238),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u104 (
		.sel (addra_pipe_0_net),
		.i0 (net_236),
		.i1 (net_240),
		.o (net_242)
	);
fifo2ram_emb_v1_AND u105 (
		.i0 (net_244),
		.i1 (net_243),
		.o (net_234)
	);
fifo2ram_emb_v1_AND u106 (
		.i0 (net_244),
		.i1 (ar[0]),
		.o (net_238)
	);
fifo2ram_emb_v1_NOT u107 (
		.i (ar[0]),
		.o (net_243)
	);
fifo2ram_emb_v1_MUX u108 (
		.sel (addra_pipe_1_net),
		.i0 (net_231),
		.i1 (net_242),
		.o (net_245)
	);
fifo2ram_emb_v1_AND u109 (
		.i0 (net_247),
		.i1 (net_246),
		.o (net_233)
	);
fifo2ram_emb_v1_AND u110 (
		.i0 (net_247),
		.i1 (ar[1]),
		.o (net_244)
	);
fifo2ram_emb_v1_NOT u111 (
		.i (ar[1]),
		.o (net_246)
	);
fifo2ram_emb_v1_MUX u112 (
		.sel (addra_pipe_2_net),
		.i0 (net_220),
		.i1 (net_245),
		.o (net_248)
	);
fifo2ram_emb_v1_AND u113 (
		.i0 (net_250),
		.i1 (net_249),
		.o (net_222)
	);
fifo2ram_emb_v1_AND u114 (
		.i0 (net_250),
		.i1 (ar[2]),
		.o (net_247)
	);
fifo2ram_emb_v1_NOT u115 (
		.i (ar[2]),
		.o (net_249)
	);
fifo2ram_emb_v1_MUX u116 (
		.sel (addra_pipe_3_net),
		.i0 (net_195),
		.i1 (net_248),
		.o (qr[1])
	);
fifo2ram_emb_v1_AND u117 (
		.i0 (cer),
		.i1 (net_252),
		.o (net_197)
	);
fifo2ram_emb_v1_AND u118 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_250)
	);
fifo2ram_emb_v1_NOT u119 (
		.i (ar[3]),
		.o (net_252)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_128 (
		.doa ({nc20161, nc20162, nc20163, nc20164, nc20165, nc20166, nc20167, nc20168, nc20169, nc20170, nc20171, nc20172, nc20173, nc20174, nc20175, nc20176, nc20177, nc20178, nc20179, nc20180, nc20181, nc20182, nc20183, nc20184, nc20185, nc20186, nc20187, nc20188, nc20189, nc20190, nc20191, nc20192, nc20193, nc20194, nc20195, nc20196, nc20197, nc20198, nc20199, nc20200, nc20201, nc20202, nc20203, nc20204, nc20205, nc20206, nc20207, nc20208, nc20209, nc20210, nc20211, nc20212, nc20213, nc20214, nc20215, nc20216, nc20217, nc20218, nc20219, nc20220, nc20221, nc20222, nc20223, net_256}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20224, nc20225, nc20226, nc20227, nc20228, nc20229, nc20230, nc20231, nc20232, nc20233, nc20234, nc20235, nc20236, nc20237, nc20238, nc20239, nc20240, nc20241, nc20242, nc20243, nc20244, nc20245, nc20246, nc20247, nc20248, nc20249, nc20250, nc20251, nc20252, nc20253, nc20254, nc20255, nc20256, nc20257, nc20258, nc20259, nc20260, nc20261, nc20262, nc20263, nc20264, nc20265, nc20266, nc20267, nc20268, nc20269, nc20270, nc20271, nc20272, nc20273, nc20274, nc20275, nc20276, nc20277, nc20278, nc20279, nc20280, nc20281, nc20282, nc20283, nc20284, nc20285, nc20286, dw[2]}),
		.dipa (),
		.dipb (),
		.cea (net_254),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_132 (
		.doa ({nc20287, nc20288, nc20289, nc20290, nc20291, nc20292, nc20293, nc20294, nc20295, nc20296, nc20297, nc20298, nc20299, nc20300, nc20301, nc20302, nc20303, nc20304, nc20305, nc20306, nc20307, nc20308, nc20309, nc20310, nc20311, nc20312, nc20313, nc20314, nc20315, nc20316, nc20317, nc20318, nc20319, nc20320, nc20321, nc20322, nc20323, nc20324, nc20325, nc20326, nc20327, nc20328, nc20329, nc20330, nc20331, nc20332, nc20333, nc20334, nc20335, nc20336, nc20337, nc20338, nc20339, nc20340, nc20341, nc20342, nc20343, nc20344, nc20345, nc20346, nc20347, nc20348, nc20349, net_260}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20350, nc20351, nc20352, nc20353, nc20354, nc20355, nc20356, nc20357, nc20358, nc20359, nc20360, nc20361, nc20362, nc20363, nc20364, nc20365, nc20366, nc20367, nc20368, nc20369, nc20370, nc20371, nc20372, nc20373, nc20374, nc20375, nc20376, nc20377, nc20378, nc20379, nc20380, nc20381, nc20382, nc20383, nc20384, nc20385, nc20386, nc20387, nc20388, nc20389, nc20390, nc20391, nc20392, nc20393, nc20394, nc20395, nc20396, nc20397, nc20398, nc20399, nc20400, nc20401, nc20402, nc20403, nc20404, nc20405, nc20406, nc20407, nc20408, nc20409, nc20410, nc20411, nc20412, dw[10]}),
		.dipa (),
		.dipb (),
		.cea (net_258),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u120 (
		.sel (addra_pipe_0_net),
		.i0 (net_256),
		.i1 (net_260),
		.o (net_262)
	);
fifo2ram_emb_v1_AND u121 (
		.i0 (net_264),
		.i1 (net_263),
		.o (net_254)
	);
fifo2ram_emb_v1_AND u122 (
		.i0 (net_264),
		.i1 (ar[0]),
		.o (net_258)
	);
fifo2ram_emb_v1_NOT u123 (
		.i (ar[0]),
		.o (net_263)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_136 (
		.doa ({nc20413, nc20414, nc20415, nc20416, nc20417, nc20418, nc20419, nc20420, nc20421, nc20422, nc20423, nc20424, nc20425, nc20426, nc20427, nc20428, nc20429, nc20430, nc20431, nc20432, nc20433, nc20434, nc20435, nc20436, nc20437, nc20438, nc20439, nc20440, nc20441, nc20442, nc20443, nc20444, nc20445, nc20446, nc20447, nc20448, nc20449, nc20450, nc20451, nc20452, nc20453, nc20454, nc20455, nc20456, nc20457, nc20458, nc20459, nc20460, nc20461, nc20462, nc20463, nc20464, nc20465, nc20466, nc20467, nc20468, nc20469, nc20470, nc20471, nc20472, nc20473, nc20474, nc20475, net_267}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20476, nc20477, nc20478, nc20479, nc20480, nc20481, nc20482, nc20483, nc20484, nc20485, nc20486, nc20487, nc20488, nc20489, nc20490, nc20491, nc20492, nc20493, nc20494, nc20495, nc20496, nc20497, nc20498, nc20499, nc20500, nc20501, nc20502, nc20503, nc20504, nc20505, nc20506, nc20507, nc20508, nc20509, nc20510, nc20511, nc20512, nc20513, nc20514, nc20515, nc20516, nc20517, nc20518, nc20519, nc20520, nc20521, nc20522, nc20523, nc20524, nc20525, nc20526, nc20527, nc20528, nc20529, nc20530, nc20531, nc20532, nc20533, nc20534, nc20535, nc20536, nc20537, nc20538, dw[18]}),
		.dipa (),
		.dipb (),
		.cea (net_265),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_140 (
		.doa ({nc20539, nc20540, nc20541, nc20542, nc20543, nc20544, nc20545, nc20546, nc20547, nc20548, nc20549, nc20550, nc20551, nc20552, nc20553, nc20554, nc20555, nc20556, nc20557, nc20558, nc20559, nc20560, nc20561, nc20562, nc20563, nc20564, nc20565, nc20566, nc20567, nc20568, nc20569, nc20570, nc20571, nc20572, nc20573, nc20574, nc20575, nc20576, nc20577, nc20578, nc20579, nc20580, nc20581, nc20582, nc20583, nc20584, nc20585, nc20586, nc20587, nc20588, nc20589, nc20590, nc20591, nc20592, nc20593, nc20594, nc20595, nc20596, nc20597, nc20598, nc20599, nc20600, nc20601, net_271}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20602, nc20603, nc20604, nc20605, nc20606, nc20607, nc20608, nc20609, nc20610, nc20611, nc20612, nc20613, nc20614, nc20615, nc20616, nc20617, nc20618, nc20619, nc20620, nc20621, nc20622, nc20623, nc20624, nc20625, nc20626, nc20627, nc20628, nc20629, nc20630, nc20631, nc20632, nc20633, nc20634, nc20635, nc20636, nc20637, nc20638, nc20639, nc20640, nc20641, nc20642, nc20643, nc20644, nc20645, nc20646, nc20647, nc20648, nc20649, nc20650, nc20651, nc20652, nc20653, nc20654, nc20655, nc20656, nc20657, nc20658, nc20659, nc20660, nc20661, nc20662, nc20663, nc20664, dw[26]}),
		.dipa (),
		.dipb (),
		.cea (net_269),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u124 (
		.sel (addra_pipe_0_net),
		.i0 (net_267),
		.i1 (net_271),
		.o (net_273)
	);
fifo2ram_emb_v1_AND u125 (
		.i0 (net_275),
		.i1 (net_274),
		.o (net_265)
	);
fifo2ram_emb_v1_AND u126 (
		.i0 (net_275),
		.i1 (ar[0]),
		.o (net_269)
	);
fifo2ram_emb_v1_NOT u127 (
		.i (ar[0]),
		.o (net_274)
	);
fifo2ram_emb_v1_MUX u128 (
		.sel (addra_pipe_1_net),
		.i0 (net_262),
		.i1 (net_273),
		.o (net_276)
	);
fifo2ram_emb_v1_AND u129 (
		.i0 (net_278),
		.i1 (net_277),
		.o (net_264)
	);
fifo2ram_emb_v1_AND u130 (
		.i0 (net_278),
		.i1 (ar[1]),
		.o (net_275)
	);
fifo2ram_emb_v1_NOT u131 (
		.i (ar[1]),
		.o (net_277)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_144 (
		.doa ({nc20665, nc20666, nc20667, nc20668, nc20669, nc20670, nc20671, nc20672, nc20673, nc20674, nc20675, nc20676, nc20677, nc20678, nc20679, nc20680, nc20681, nc20682, nc20683, nc20684, nc20685, nc20686, nc20687, nc20688, nc20689, nc20690, nc20691, nc20692, nc20693, nc20694, nc20695, nc20696, nc20697, nc20698, nc20699, nc20700, nc20701, nc20702, nc20703, nc20704, nc20705, nc20706, nc20707, nc20708, nc20709, nc20710, nc20711, nc20712, nc20713, nc20714, nc20715, nc20716, nc20717, nc20718, nc20719, nc20720, nc20721, nc20722, nc20723, nc20724, nc20725, nc20726, nc20727, net_281}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20728, nc20729, nc20730, nc20731, nc20732, nc20733, nc20734, nc20735, nc20736, nc20737, nc20738, nc20739, nc20740, nc20741, nc20742, nc20743, nc20744, nc20745, nc20746, nc20747, nc20748, nc20749, nc20750, nc20751, nc20752, nc20753, nc20754, nc20755, nc20756, nc20757, nc20758, nc20759, nc20760, nc20761, nc20762, nc20763, nc20764, nc20765, nc20766, nc20767, nc20768, nc20769, nc20770, nc20771, nc20772, nc20773, nc20774, nc20775, nc20776, nc20777, nc20778, nc20779, nc20780, nc20781, nc20782, nc20783, nc20784, nc20785, nc20786, nc20787, nc20788, nc20789, nc20790, dw[34]}),
		.dipa (),
		.dipb (),
		.cea (net_279),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_148 (
		.doa ({nc20791, nc20792, nc20793, nc20794, nc20795, nc20796, nc20797, nc20798, nc20799, nc20800, nc20801, nc20802, nc20803, nc20804, nc20805, nc20806, nc20807, nc20808, nc20809, nc20810, nc20811, nc20812, nc20813, nc20814, nc20815, nc20816, nc20817, nc20818, nc20819, nc20820, nc20821, nc20822, nc20823, nc20824, nc20825, nc20826, nc20827, nc20828, nc20829, nc20830, nc20831, nc20832, nc20833, nc20834, nc20835, nc20836, nc20837, nc20838, nc20839, nc20840, nc20841, nc20842, nc20843, nc20844, nc20845, nc20846, nc20847, nc20848, nc20849, nc20850, nc20851, nc20852, nc20853, net_285}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20854, nc20855, nc20856, nc20857, nc20858, nc20859, nc20860, nc20861, nc20862, nc20863, nc20864, nc20865, nc20866, nc20867, nc20868, nc20869, nc20870, nc20871, nc20872, nc20873, nc20874, nc20875, nc20876, nc20877, nc20878, nc20879, nc20880, nc20881, nc20882, nc20883, nc20884, nc20885, nc20886, nc20887, nc20888, nc20889, nc20890, nc20891, nc20892, nc20893, nc20894, nc20895, nc20896, nc20897, nc20898, nc20899, nc20900, nc20901, nc20902, nc20903, nc20904, nc20905, nc20906, nc20907, nc20908, nc20909, nc20910, nc20911, nc20912, nc20913, nc20914, nc20915, nc20916, dw[42]}),
		.dipa (),
		.dipb (),
		.cea (net_283),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u132 (
		.sel (addra_pipe_0_net),
		.i0 (net_281),
		.i1 (net_285),
		.o (net_287)
	);
fifo2ram_emb_v1_AND u133 (
		.i0 (net_289),
		.i1 (net_288),
		.o (net_279)
	);
fifo2ram_emb_v1_AND u134 (
		.i0 (net_289),
		.i1 (ar[0]),
		.o (net_283)
	);
fifo2ram_emb_v1_NOT u135 (
		.i (ar[0]),
		.o (net_288)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_152 (
		.doa ({nc20917, nc20918, nc20919, nc20920, nc20921, nc20922, nc20923, nc20924, nc20925, nc20926, nc20927, nc20928, nc20929, nc20930, nc20931, nc20932, nc20933, nc20934, nc20935, nc20936, nc20937, nc20938, nc20939, nc20940, nc20941, nc20942, nc20943, nc20944, nc20945, nc20946, nc20947, nc20948, nc20949, nc20950, nc20951, nc20952, nc20953, nc20954, nc20955, nc20956, nc20957, nc20958, nc20959, nc20960, nc20961, nc20962, nc20963, nc20964, nc20965, nc20966, nc20967, nc20968, nc20969, nc20970, nc20971, nc20972, nc20973, nc20974, nc20975, nc20976, nc20977, nc20978, nc20979, net_292}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc20980, nc20981, nc20982, nc20983, nc20984, nc20985, nc20986, nc20987, nc20988, nc20989, nc20990, nc20991, nc20992, nc20993, nc20994, nc20995, nc20996, nc20997, nc20998, nc20999, nc21000, nc21001, nc21002, nc21003, nc21004, nc21005, nc21006, nc21007, nc21008, nc21009, nc21010, nc21011, nc21012, nc21013, nc21014, nc21015, nc21016, nc21017, nc21018, nc21019, nc21020, nc21021, nc21022, nc21023, nc21024, nc21025, nc21026, nc21027, nc21028, nc21029, nc21030, nc21031, nc21032, nc21033, nc21034, nc21035, nc21036, nc21037, nc21038, nc21039, nc21040, nc21041, nc21042, dw[50]}),
		.dipa (),
		.dipb (),
		.cea (net_290),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_156 (
		.doa ({nc21043, nc21044, nc21045, nc21046, nc21047, nc21048, nc21049, nc21050, nc21051, nc21052, nc21053, nc21054, nc21055, nc21056, nc21057, nc21058, nc21059, nc21060, nc21061, nc21062, nc21063, nc21064, nc21065, nc21066, nc21067, nc21068, nc21069, nc21070, nc21071, nc21072, nc21073, nc21074, nc21075, nc21076, nc21077, nc21078, nc21079, nc21080, nc21081, nc21082, nc21083, nc21084, nc21085, nc21086, nc21087, nc21088, nc21089, nc21090, nc21091, nc21092, nc21093, nc21094, nc21095, nc21096, nc21097, nc21098, nc21099, nc21100, nc21101, nc21102, nc21103, nc21104, nc21105, net_296}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21106, nc21107, nc21108, nc21109, nc21110, nc21111, nc21112, nc21113, nc21114, nc21115, nc21116, nc21117, nc21118, nc21119, nc21120, nc21121, nc21122, nc21123, nc21124, nc21125, nc21126, nc21127, nc21128, nc21129, nc21130, nc21131, nc21132, nc21133, nc21134, nc21135, nc21136, nc21137, nc21138, nc21139, nc21140, nc21141, nc21142, nc21143, nc21144, nc21145, nc21146, nc21147, nc21148, nc21149, nc21150, nc21151, nc21152, nc21153, nc21154, nc21155, nc21156, nc21157, nc21158, nc21159, nc21160, nc21161, nc21162, nc21163, nc21164, nc21165, nc21166, nc21167, nc21168, dw[58]}),
		.dipa (),
		.dipb (),
		.cea (net_294),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u136 (
		.sel (addra_pipe_0_net),
		.i0 (net_292),
		.i1 (net_296),
		.o (net_298)
	);
fifo2ram_emb_v1_AND u137 (
		.i0 (net_300),
		.i1 (net_299),
		.o (net_290)
	);
fifo2ram_emb_v1_AND u138 (
		.i0 (net_300),
		.i1 (ar[0]),
		.o (net_294)
	);
fifo2ram_emb_v1_NOT u139 (
		.i (ar[0]),
		.o (net_299)
	);
fifo2ram_emb_v1_MUX u140 (
		.sel (addra_pipe_1_net),
		.i0 (net_287),
		.i1 (net_298),
		.o (net_301)
	);
fifo2ram_emb_v1_AND u141 (
		.i0 (net_303),
		.i1 (net_302),
		.o (net_289)
	);
fifo2ram_emb_v1_AND u142 (
		.i0 (net_303),
		.i1 (ar[1]),
		.o (net_300)
	);
fifo2ram_emb_v1_NOT u143 (
		.i (ar[1]),
		.o (net_302)
	);
fifo2ram_emb_v1_MUX u144 (
		.sel (addra_pipe_2_net),
		.i0 (net_276),
		.i1 (net_301),
		.o (net_304)
	);
fifo2ram_emb_v1_AND u145 (
		.i0 (net_306),
		.i1 (net_305),
		.o (net_278)
	);
fifo2ram_emb_v1_AND u146 (
		.i0 (net_306),
		.i1 (ar[2]),
		.o (net_303)
	);
fifo2ram_emb_v1_NOT u147 (
		.i (ar[2]),
		.o (net_305)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_160 (
		.doa ({nc21169, nc21170, nc21171, nc21172, nc21173, nc21174, nc21175, nc21176, nc21177, nc21178, nc21179, nc21180, nc21181, nc21182, nc21183, nc21184, nc21185, nc21186, nc21187, nc21188, nc21189, nc21190, nc21191, nc21192, nc21193, nc21194, nc21195, nc21196, nc21197, nc21198, nc21199, nc21200, nc21201, nc21202, nc21203, nc21204, nc21205, nc21206, nc21207, nc21208, nc21209, nc21210, nc21211, nc21212, nc21213, nc21214, nc21215, nc21216, nc21217, nc21218, nc21219, nc21220, nc21221, nc21222, nc21223, nc21224, nc21225, nc21226, nc21227, nc21228, nc21229, nc21230, nc21231, net_309}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21232, nc21233, nc21234, nc21235, nc21236, nc21237, nc21238, nc21239, nc21240, nc21241, nc21242, nc21243, nc21244, nc21245, nc21246, nc21247, nc21248, nc21249, nc21250, nc21251, nc21252, nc21253, nc21254, nc21255, nc21256, nc21257, nc21258, nc21259, nc21260, nc21261, nc21262, nc21263, nc21264, nc21265, nc21266, nc21267, nc21268, nc21269, nc21270, nc21271, nc21272, nc21273, nc21274, nc21275, nc21276, nc21277, nc21278, nc21279, nc21280, nc21281, nc21282, nc21283, nc21284, nc21285, nc21286, nc21287, nc21288, nc21289, nc21290, nc21291, nc21292, nc21293, nc21294, dw[66]}),
		.dipa (),
		.dipb (),
		.cea (net_307),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_164 (
		.doa ({nc21295, nc21296, nc21297, nc21298, nc21299, nc21300, nc21301, nc21302, nc21303, nc21304, nc21305, nc21306, nc21307, nc21308, nc21309, nc21310, nc21311, nc21312, nc21313, nc21314, nc21315, nc21316, nc21317, nc21318, nc21319, nc21320, nc21321, nc21322, nc21323, nc21324, nc21325, nc21326, nc21327, nc21328, nc21329, nc21330, nc21331, nc21332, nc21333, nc21334, nc21335, nc21336, nc21337, nc21338, nc21339, nc21340, nc21341, nc21342, nc21343, nc21344, nc21345, nc21346, nc21347, nc21348, nc21349, nc21350, nc21351, nc21352, nc21353, nc21354, nc21355, nc21356, nc21357, net_313}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21358, nc21359, nc21360, nc21361, nc21362, nc21363, nc21364, nc21365, nc21366, nc21367, nc21368, nc21369, nc21370, nc21371, nc21372, nc21373, nc21374, nc21375, nc21376, nc21377, nc21378, nc21379, nc21380, nc21381, nc21382, nc21383, nc21384, nc21385, nc21386, nc21387, nc21388, nc21389, nc21390, nc21391, nc21392, nc21393, nc21394, nc21395, nc21396, nc21397, nc21398, nc21399, nc21400, nc21401, nc21402, nc21403, nc21404, nc21405, nc21406, nc21407, nc21408, nc21409, nc21410, nc21411, nc21412, nc21413, nc21414, nc21415, nc21416, nc21417, nc21418, nc21419, nc21420, dw[74]}),
		.dipa (),
		.dipb (),
		.cea (net_311),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u148 (
		.sel (addra_pipe_0_net),
		.i0 (net_309),
		.i1 (net_313),
		.o (net_315)
	);
fifo2ram_emb_v1_AND u149 (
		.i0 (net_317),
		.i1 (net_316),
		.o (net_307)
	);
fifo2ram_emb_v1_AND u150 (
		.i0 (net_317),
		.i1 (ar[0]),
		.o (net_311)
	);
fifo2ram_emb_v1_NOT u151 (
		.i (ar[0]),
		.o (net_316)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_168 (
		.doa ({nc21421, nc21422, nc21423, nc21424, nc21425, nc21426, nc21427, nc21428, nc21429, nc21430, nc21431, nc21432, nc21433, nc21434, nc21435, nc21436, nc21437, nc21438, nc21439, nc21440, nc21441, nc21442, nc21443, nc21444, nc21445, nc21446, nc21447, nc21448, nc21449, nc21450, nc21451, nc21452, nc21453, nc21454, nc21455, nc21456, nc21457, nc21458, nc21459, nc21460, nc21461, nc21462, nc21463, nc21464, nc21465, nc21466, nc21467, nc21468, nc21469, nc21470, nc21471, nc21472, nc21473, nc21474, nc21475, nc21476, nc21477, nc21478, nc21479, nc21480, nc21481, nc21482, nc21483, net_320}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21484, nc21485, nc21486, nc21487, nc21488, nc21489, nc21490, nc21491, nc21492, nc21493, nc21494, nc21495, nc21496, nc21497, nc21498, nc21499, nc21500, nc21501, nc21502, nc21503, nc21504, nc21505, nc21506, nc21507, nc21508, nc21509, nc21510, nc21511, nc21512, nc21513, nc21514, nc21515, nc21516, nc21517, nc21518, nc21519, nc21520, nc21521, nc21522, nc21523, nc21524, nc21525, nc21526, nc21527, nc21528, nc21529, nc21530, nc21531, nc21532, nc21533, nc21534, nc21535, nc21536, nc21537, nc21538, nc21539, nc21540, nc21541, nc21542, nc21543, nc21544, nc21545, nc21546, dw[82]}),
		.dipa (),
		.dipb (),
		.cea (net_318),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_172 (
		.doa ({nc21547, nc21548, nc21549, nc21550, nc21551, nc21552, nc21553, nc21554, nc21555, nc21556, nc21557, nc21558, nc21559, nc21560, nc21561, nc21562, nc21563, nc21564, nc21565, nc21566, nc21567, nc21568, nc21569, nc21570, nc21571, nc21572, nc21573, nc21574, nc21575, nc21576, nc21577, nc21578, nc21579, nc21580, nc21581, nc21582, nc21583, nc21584, nc21585, nc21586, nc21587, nc21588, nc21589, nc21590, nc21591, nc21592, nc21593, nc21594, nc21595, nc21596, nc21597, nc21598, nc21599, nc21600, nc21601, nc21602, nc21603, nc21604, nc21605, nc21606, nc21607, nc21608, nc21609, net_324}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21610, nc21611, nc21612, nc21613, nc21614, nc21615, nc21616, nc21617, nc21618, nc21619, nc21620, nc21621, nc21622, nc21623, nc21624, nc21625, nc21626, nc21627, nc21628, nc21629, nc21630, nc21631, nc21632, nc21633, nc21634, nc21635, nc21636, nc21637, nc21638, nc21639, nc21640, nc21641, nc21642, nc21643, nc21644, nc21645, nc21646, nc21647, nc21648, nc21649, nc21650, nc21651, nc21652, nc21653, nc21654, nc21655, nc21656, nc21657, nc21658, nc21659, nc21660, nc21661, nc21662, nc21663, nc21664, nc21665, nc21666, nc21667, nc21668, nc21669, nc21670, nc21671, nc21672, dw[90]}),
		.dipa (),
		.dipb (),
		.cea (net_322),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u152 (
		.sel (addra_pipe_0_net),
		.i0 (net_320),
		.i1 (net_324),
		.o (net_326)
	);
fifo2ram_emb_v1_AND u153 (
		.i0 (net_328),
		.i1 (net_327),
		.o (net_318)
	);
fifo2ram_emb_v1_AND u154 (
		.i0 (net_328),
		.i1 (ar[0]),
		.o (net_322)
	);
fifo2ram_emb_v1_NOT u155 (
		.i (ar[0]),
		.o (net_327)
	);
fifo2ram_emb_v1_MUX u156 (
		.sel (addra_pipe_1_net),
		.i0 (net_315),
		.i1 (net_326),
		.o (net_329)
	);
fifo2ram_emb_v1_AND u157 (
		.i0 (net_331),
		.i1 (net_330),
		.o (net_317)
	);
fifo2ram_emb_v1_AND u158 (
		.i0 (net_331),
		.i1 (ar[1]),
		.o (net_328)
	);
fifo2ram_emb_v1_NOT u159 (
		.i (ar[1]),
		.o (net_330)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_176 (
		.doa ({nc21673, nc21674, nc21675, nc21676, nc21677, nc21678, nc21679, nc21680, nc21681, nc21682, nc21683, nc21684, nc21685, nc21686, nc21687, nc21688, nc21689, nc21690, nc21691, nc21692, nc21693, nc21694, nc21695, nc21696, nc21697, nc21698, nc21699, nc21700, nc21701, nc21702, nc21703, nc21704, nc21705, nc21706, nc21707, nc21708, nc21709, nc21710, nc21711, nc21712, nc21713, nc21714, nc21715, nc21716, nc21717, nc21718, nc21719, nc21720, nc21721, nc21722, nc21723, nc21724, nc21725, nc21726, nc21727, nc21728, nc21729, nc21730, nc21731, nc21732, nc21733, nc21734, nc21735, net_334}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21736, nc21737, nc21738, nc21739, nc21740, nc21741, nc21742, nc21743, nc21744, nc21745, nc21746, nc21747, nc21748, nc21749, nc21750, nc21751, nc21752, nc21753, nc21754, nc21755, nc21756, nc21757, nc21758, nc21759, nc21760, nc21761, nc21762, nc21763, nc21764, nc21765, nc21766, nc21767, nc21768, nc21769, nc21770, nc21771, nc21772, nc21773, nc21774, nc21775, nc21776, nc21777, nc21778, nc21779, nc21780, nc21781, nc21782, nc21783, nc21784, nc21785, nc21786, nc21787, nc21788, nc21789, nc21790, nc21791, nc21792, nc21793, nc21794, nc21795, nc21796, nc21797, nc21798, dw[98]}),
		.dipa (),
		.dipb (),
		.cea (net_332),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_180 (
		.doa ({nc21799, nc21800, nc21801, nc21802, nc21803, nc21804, nc21805, nc21806, nc21807, nc21808, nc21809, nc21810, nc21811, nc21812, nc21813, nc21814, nc21815, nc21816, nc21817, nc21818, nc21819, nc21820, nc21821, nc21822, nc21823, nc21824, nc21825, nc21826, nc21827, nc21828, nc21829, nc21830, nc21831, nc21832, nc21833, nc21834, nc21835, nc21836, nc21837, nc21838, nc21839, nc21840, nc21841, nc21842, nc21843, nc21844, nc21845, nc21846, nc21847, nc21848, nc21849, nc21850, nc21851, nc21852, nc21853, nc21854, nc21855, nc21856, nc21857, nc21858, nc21859, nc21860, nc21861, net_338}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21862, nc21863, nc21864, nc21865, nc21866, nc21867, nc21868, nc21869, nc21870, nc21871, nc21872, nc21873, nc21874, nc21875, nc21876, nc21877, nc21878, nc21879, nc21880, nc21881, nc21882, nc21883, nc21884, nc21885, nc21886, nc21887, nc21888, nc21889, nc21890, nc21891, nc21892, nc21893, nc21894, nc21895, nc21896, nc21897, nc21898, nc21899, nc21900, nc21901, nc21902, nc21903, nc21904, nc21905, nc21906, nc21907, nc21908, nc21909, nc21910, nc21911, nc21912, nc21913, nc21914, nc21915, nc21916, nc21917, nc21918, nc21919, nc21920, nc21921, nc21922, nc21923, nc21924, dw[106]}),
		.dipa (),
		.dipb (),
		.cea (net_336),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u160 (
		.sel (addra_pipe_0_net),
		.i0 (net_334),
		.i1 (net_338),
		.o (net_340)
	);
fifo2ram_emb_v1_AND u161 (
		.i0 (net_342),
		.i1 (net_341),
		.o (net_332)
	);
fifo2ram_emb_v1_AND u162 (
		.i0 (net_342),
		.i1 (ar[0]),
		.o (net_336)
	);
fifo2ram_emb_v1_NOT u163 (
		.i (ar[0]),
		.o (net_341)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_184 (
		.doa ({nc21925, nc21926, nc21927, nc21928, nc21929, nc21930, nc21931, nc21932, nc21933, nc21934, nc21935, nc21936, nc21937, nc21938, nc21939, nc21940, nc21941, nc21942, nc21943, nc21944, nc21945, nc21946, nc21947, nc21948, nc21949, nc21950, nc21951, nc21952, nc21953, nc21954, nc21955, nc21956, nc21957, nc21958, nc21959, nc21960, nc21961, nc21962, nc21963, nc21964, nc21965, nc21966, nc21967, nc21968, nc21969, nc21970, nc21971, nc21972, nc21973, nc21974, nc21975, nc21976, nc21977, nc21978, nc21979, nc21980, nc21981, nc21982, nc21983, nc21984, nc21985, nc21986, nc21987, net_345}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc21988, nc21989, nc21990, nc21991, nc21992, nc21993, nc21994, nc21995, nc21996, nc21997, nc21998, nc21999, nc22000, nc22001, nc22002, nc22003, nc22004, nc22005, nc22006, nc22007, nc22008, nc22009, nc22010, nc22011, nc22012, nc22013, nc22014, nc22015, nc22016, nc22017, nc22018, nc22019, nc22020, nc22021, nc22022, nc22023, nc22024, nc22025, nc22026, nc22027, nc22028, nc22029, nc22030, nc22031, nc22032, nc22033, nc22034, nc22035, nc22036, nc22037, nc22038, nc22039, nc22040, nc22041, nc22042, nc22043, nc22044, nc22045, nc22046, nc22047, nc22048, nc22049, nc22050, dw[114]}),
		.dipa (),
		.dipb (),
		.cea (net_343),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_188 (
		.doa ({nc22051, nc22052, nc22053, nc22054, nc22055, nc22056, nc22057, nc22058, nc22059, nc22060, nc22061, nc22062, nc22063, nc22064, nc22065, nc22066, nc22067, nc22068, nc22069, nc22070, nc22071, nc22072, nc22073, nc22074, nc22075, nc22076, nc22077, nc22078, nc22079, nc22080, nc22081, nc22082, nc22083, nc22084, nc22085, nc22086, nc22087, nc22088, nc22089, nc22090, nc22091, nc22092, nc22093, nc22094, nc22095, nc22096, nc22097, nc22098, nc22099, nc22100, nc22101, nc22102, nc22103, nc22104, nc22105, nc22106, nc22107, nc22108, nc22109, nc22110, nc22111, nc22112, nc22113, net_349}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22114, nc22115, nc22116, nc22117, nc22118, nc22119, nc22120, nc22121, nc22122, nc22123, nc22124, nc22125, nc22126, nc22127, nc22128, nc22129, nc22130, nc22131, nc22132, nc22133, nc22134, nc22135, nc22136, nc22137, nc22138, nc22139, nc22140, nc22141, nc22142, nc22143, nc22144, nc22145, nc22146, nc22147, nc22148, nc22149, nc22150, nc22151, nc22152, nc22153, nc22154, nc22155, nc22156, nc22157, nc22158, nc22159, nc22160, nc22161, nc22162, nc22163, nc22164, nc22165, nc22166, nc22167, nc22168, nc22169, nc22170, nc22171, nc22172, nc22173, nc22174, nc22175, nc22176, dw[122]}),
		.dipa (),
		.dipb (),
		.cea (net_347),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u164 (
		.sel (addra_pipe_0_net),
		.i0 (net_345),
		.i1 (net_349),
		.o (net_351)
	);
fifo2ram_emb_v1_AND u165 (
		.i0 (net_353),
		.i1 (net_352),
		.o (net_343)
	);
fifo2ram_emb_v1_AND u166 (
		.i0 (net_353),
		.i1 (ar[0]),
		.o (net_347)
	);
fifo2ram_emb_v1_NOT u167 (
		.i (ar[0]),
		.o (net_352)
	);
fifo2ram_emb_v1_MUX u168 (
		.sel (addra_pipe_1_net),
		.i0 (net_340),
		.i1 (net_351),
		.o (net_354)
	);
fifo2ram_emb_v1_AND u169 (
		.i0 (net_356),
		.i1 (net_355),
		.o (net_342)
	);
fifo2ram_emb_v1_AND u170 (
		.i0 (net_356),
		.i1 (ar[1]),
		.o (net_353)
	);
fifo2ram_emb_v1_NOT u171 (
		.i (ar[1]),
		.o (net_355)
	);
fifo2ram_emb_v1_MUX u172 (
		.sel (addra_pipe_2_net),
		.i0 (net_329),
		.i1 (net_354),
		.o (net_357)
	);
fifo2ram_emb_v1_AND u173 (
		.i0 (net_359),
		.i1 (net_358),
		.o (net_331)
	);
fifo2ram_emb_v1_AND u174 (
		.i0 (net_359),
		.i1 (ar[2]),
		.o (net_356)
	);
fifo2ram_emb_v1_NOT u175 (
		.i (ar[2]),
		.o (net_358)
	);
fifo2ram_emb_v1_MUX u176 (
		.sel (addra_pipe_3_net),
		.i0 (net_304),
		.i1 (net_357),
		.o (qr[2])
	);
fifo2ram_emb_v1_AND u177 (
		.i0 (cer),
		.i1 (net_361),
		.o (net_306)
	);
fifo2ram_emb_v1_AND u178 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_359)
	);
fifo2ram_emb_v1_NOT u179 (
		.i (ar[3]),
		.o (net_361)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_192 (
		.doa ({nc22177, nc22178, nc22179, nc22180, nc22181, nc22182, nc22183, nc22184, nc22185, nc22186, nc22187, nc22188, nc22189, nc22190, nc22191, nc22192, nc22193, nc22194, nc22195, nc22196, nc22197, nc22198, nc22199, nc22200, nc22201, nc22202, nc22203, nc22204, nc22205, nc22206, nc22207, nc22208, nc22209, nc22210, nc22211, nc22212, nc22213, nc22214, nc22215, nc22216, nc22217, nc22218, nc22219, nc22220, nc22221, nc22222, nc22223, nc22224, nc22225, nc22226, nc22227, nc22228, nc22229, nc22230, nc22231, nc22232, nc22233, nc22234, nc22235, nc22236, nc22237, nc22238, nc22239, net_365}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22240, nc22241, nc22242, nc22243, nc22244, nc22245, nc22246, nc22247, nc22248, nc22249, nc22250, nc22251, nc22252, nc22253, nc22254, nc22255, nc22256, nc22257, nc22258, nc22259, nc22260, nc22261, nc22262, nc22263, nc22264, nc22265, nc22266, nc22267, nc22268, nc22269, nc22270, nc22271, nc22272, nc22273, nc22274, nc22275, nc22276, nc22277, nc22278, nc22279, nc22280, nc22281, nc22282, nc22283, nc22284, nc22285, nc22286, nc22287, nc22288, nc22289, nc22290, nc22291, nc22292, nc22293, nc22294, nc22295, nc22296, nc22297, nc22298, nc22299, nc22300, nc22301, nc22302, dw[3]}),
		.dipa (),
		.dipb (),
		.cea (net_363),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_196 (
		.doa ({nc22303, nc22304, nc22305, nc22306, nc22307, nc22308, nc22309, nc22310, nc22311, nc22312, nc22313, nc22314, nc22315, nc22316, nc22317, nc22318, nc22319, nc22320, nc22321, nc22322, nc22323, nc22324, nc22325, nc22326, nc22327, nc22328, nc22329, nc22330, nc22331, nc22332, nc22333, nc22334, nc22335, nc22336, nc22337, nc22338, nc22339, nc22340, nc22341, nc22342, nc22343, nc22344, nc22345, nc22346, nc22347, nc22348, nc22349, nc22350, nc22351, nc22352, nc22353, nc22354, nc22355, nc22356, nc22357, nc22358, nc22359, nc22360, nc22361, nc22362, nc22363, nc22364, nc22365, net_369}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22366, nc22367, nc22368, nc22369, nc22370, nc22371, nc22372, nc22373, nc22374, nc22375, nc22376, nc22377, nc22378, nc22379, nc22380, nc22381, nc22382, nc22383, nc22384, nc22385, nc22386, nc22387, nc22388, nc22389, nc22390, nc22391, nc22392, nc22393, nc22394, nc22395, nc22396, nc22397, nc22398, nc22399, nc22400, nc22401, nc22402, nc22403, nc22404, nc22405, nc22406, nc22407, nc22408, nc22409, nc22410, nc22411, nc22412, nc22413, nc22414, nc22415, nc22416, nc22417, nc22418, nc22419, nc22420, nc22421, nc22422, nc22423, nc22424, nc22425, nc22426, nc22427, nc22428, dw[11]}),
		.dipa (),
		.dipb (),
		.cea (net_367),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u180 (
		.sel (addra_pipe_0_net),
		.i0 (net_365),
		.i1 (net_369),
		.o (net_371)
	);
fifo2ram_emb_v1_AND u181 (
		.i0 (net_373),
		.i1 (net_372),
		.o (net_363)
	);
fifo2ram_emb_v1_AND u182 (
		.i0 (net_373),
		.i1 (ar[0]),
		.o (net_367)
	);
fifo2ram_emb_v1_NOT u183 (
		.i (ar[0]),
		.o (net_372)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_200 (
		.doa ({nc22429, nc22430, nc22431, nc22432, nc22433, nc22434, nc22435, nc22436, nc22437, nc22438, nc22439, nc22440, nc22441, nc22442, nc22443, nc22444, nc22445, nc22446, nc22447, nc22448, nc22449, nc22450, nc22451, nc22452, nc22453, nc22454, nc22455, nc22456, nc22457, nc22458, nc22459, nc22460, nc22461, nc22462, nc22463, nc22464, nc22465, nc22466, nc22467, nc22468, nc22469, nc22470, nc22471, nc22472, nc22473, nc22474, nc22475, nc22476, nc22477, nc22478, nc22479, nc22480, nc22481, nc22482, nc22483, nc22484, nc22485, nc22486, nc22487, nc22488, nc22489, nc22490, nc22491, net_376}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22492, nc22493, nc22494, nc22495, nc22496, nc22497, nc22498, nc22499, nc22500, nc22501, nc22502, nc22503, nc22504, nc22505, nc22506, nc22507, nc22508, nc22509, nc22510, nc22511, nc22512, nc22513, nc22514, nc22515, nc22516, nc22517, nc22518, nc22519, nc22520, nc22521, nc22522, nc22523, nc22524, nc22525, nc22526, nc22527, nc22528, nc22529, nc22530, nc22531, nc22532, nc22533, nc22534, nc22535, nc22536, nc22537, nc22538, nc22539, nc22540, nc22541, nc22542, nc22543, nc22544, nc22545, nc22546, nc22547, nc22548, nc22549, nc22550, nc22551, nc22552, nc22553, nc22554, dw[19]}),
		.dipa (),
		.dipb (),
		.cea (net_374),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_204 (
		.doa ({nc22555, nc22556, nc22557, nc22558, nc22559, nc22560, nc22561, nc22562, nc22563, nc22564, nc22565, nc22566, nc22567, nc22568, nc22569, nc22570, nc22571, nc22572, nc22573, nc22574, nc22575, nc22576, nc22577, nc22578, nc22579, nc22580, nc22581, nc22582, nc22583, nc22584, nc22585, nc22586, nc22587, nc22588, nc22589, nc22590, nc22591, nc22592, nc22593, nc22594, nc22595, nc22596, nc22597, nc22598, nc22599, nc22600, nc22601, nc22602, nc22603, nc22604, nc22605, nc22606, nc22607, nc22608, nc22609, nc22610, nc22611, nc22612, nc22613, nc22614, nc22615, nc22616, nc22617, net_380}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22618, nc22619, nc22620, nc22621, nc22622, nc22623, nc22624, nc22625, nc22626, nc22627, nc22628, nc22629, nc22630, nc22631, nc22632, nc22633, nc22634, nc22635, nc22636, nc22637, nc22638, nc22639, nc22640, nc22641, nc22642, nc22643, nc22644, nc22645, nc22646, nc22647, nc22648, nc22649, nc22650, nc22651, nc22652, nc22653, nc22654, nc22655, nc22656, nc22657, nc22658, nc22659, nc22660, nc22661, nc22662, nc22663, nc22664, nc22665, nc22666, nc22667, nc22668, nc22669, nc22670, nc22671, nc22672, nc22673, nc22674, nc22675, nc22676, nc22677, nc22678, nc22679, nc22680, dw[27]}),
		.dipa (),
		.dipb (),
		.cea (net_378),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u184 (
		.sel (addra_pipe_0_net),
		.i0 (net_376),
		.i1 (net_380),
		.o (net_382)
	);
fifo2ram_emb_v1_AND u185 (
		.i0 (net_384),
		.i1 (net_383),
		.o (net_374)
	);
fifo2ram_emb_v1_AND u186 (
		.i0 (net_384),
		.i1 (ar[0]),
		.o (net_378)
	);
fifo2ram_emb_v1_NOT u187 (
		.i (ar[0]),
		.o (net_383)
	);
fifo2ram_emb_v1_MUX u188 (
		.sel (addra_pipe_1_net),
		.i0 (net_371),
		.i1 (net_382),
		.o (net_385)
	);
fifo2ram_emb_v1_AND u189 (
		.i0 (net_387),
		.i1 (net_386),
		.o (net_373)
	);
fifo2ram_emb_v1_AND u190 (
		.i0 (net_387),
		.i1 (ar[1]),
		.o (net_384)
	);
fifo2ram_emb_v1_NOT u191 (
		.i (ar[1]),
		.o (net_386)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_208 (
		.doa ({nc22681, nc22682, nc22683, nc22684, nc22685, nc22686, nc22687, nc22688, nc22689, nc22690, nc22691, nc22692, nc22693, nc22694, nc22695, nc22696, nc22697, nc22698, nc22699, nc22700, nc22701, nc22702, nc22703, nc22704, nc22705, nc22706, nc22707, nc22708, nc22709, nc22710, nc22711, nc22712, nc22713, nc22714, nc22715, nc22716, nc22717, nc22718, nc22719, nc22720, nc22721, nc22722, nc22723, nc22724, nc22725, nc22726, nc22727, nc22728, nc22729, nc22730, nc22731, nc22732, nc22733, nc22734, nc22735, nc22736, nc22737, nc22738, nc22739, nc22740, nc22741, nc22742, nc22743, net_390}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22744, nc22745, nc22746, nc22747, nc22748, nc22749, nc22750, nc22751, nc22752, nc22753, nc22754, nc22755, nc22756, nc22757, nc22758, nc22759, nc22760, nc22761, nc22762, nc22763, nc22764, nc22765, nc22766, nc22767, nc22768, nc22769, nc22770, nc22771, nc22772, nc22773, nc22774, nc22775, nc22776, nc22777, nc22778, nc22779, nc22780, nc22781, nc22782, nc22783, nc22784, nc22785, nc22786, nc22787, nc22788, nc22789, nc22790, nc22791, nc22792, nc22793, nc22794, nc22795, nc22796, nc22797, nc22798, nc22799, nc22800, nc22801, nc22802, nc22803, nc22804, nc22805, nc22806, dw[35]}),
		.dipa (),
		.dipb (),
		.cea (net_388),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_212 (
		.doa ({nc22807, nc22808, nc22809, nc22810, nc22811, nc22812, nc22813, nc22814, nc22815, nc22816, nc22817, nc22818, nc22819, nc22820, nc22821, nc22822, nc22823, nc22824, nc22825, nc22826, nc22827, nc22828, nc22829, nc22830, nc22831, nc22832, nc22833, nc22834, nc22835, nc22836, nc22837, nc22838, nc22839, nc22840, nc22841, nc22842, nc22843, nc22844, nc22845, nc22846, nc22847, nc22848, nc22849, nc22850, nc22851, nc22852, nc22853, nc22854, nc22855, nc22856, nc22857, nc22858, nc22859, nc22860, nc22861, nc22862, nc22863, nc22864, nc22865, nc22866, nc22867, nc22868, nc22869, net_394}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22870, nc22871, nc22872, nc22873, nc22874, nc22875, nc22876, nc22877, nc22878, nc22879, nc22880, nc22881, nc22882, nc22883, nc22884, nc22885, nc22886, nc22887, nc22888, nc22889, nc22890, nc22891, nc22892, nc22893, nc22894, nc22895, nc22896, nc22897, nc22898, nc22899, nc22900, nc22901, nc22902, nc22903, nc22904, nc22905, nc22906, nc22907, nc22908, nc22909, nc22910, nc22911, nc22912, nc22913, nc22914, nc22915, nc22916, nc22917, nc22918, nc22919, nc22920, nc22921, nc22922, nc22923, nc22924, nc22925, nc22926, nc22927, nc22928, nc22929, nc22930, nc22931, nc22932, dw[43]}),
		.dipa (),
		.dipb (),
		.cea (net_392),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u192 (
		.sel (addra_pipe_0_net),
		.i0 (net_390),
		.i1 (net_394),
		.o (net_396)
	);
fifo2ram_emb_v1_AND u193 (
		.i0 (net_398),
		.i1 (net_397),
		.o (net_388)
	);
fifo2ram_emb_v1_AND u194 (
		.i0 (net_398),
		.i1 (ar[0]),
		.o (net_392)
	);
fifo2ram_emb_v1_NOT u195 (
		.i (ar[0]),
		.o (net_397)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_216 (
		.doa ({nc22933, nc22934, nc22935, nc22936, nc22937, nc22938, nc22939, nc22940, nc22941, nc22942, nc22943, nc22944, nc22945, nc22946, nc22947, nc22948, nc22949, nc22950, nc22951, nc22952, nc22953, nc22954, nc22955, nc22956, nc22957, nc22958, nc22959, nc22960, nc22961, nc22962, nc22963, nc22964, nc22965, nc22966, nc22967, nc22968, nc22969, nc22970, nc22971, nc22972, nc22973, nc22974, nc22975, nc22976, nc22977, nc22978, nc22979, nc22980, nc22981, nc22982, nc22983, nc22984, nc22985, nc22986, nc22987, nc22988, nc22989, nc22990, nc22991, nc22992, nc22993, nc22994, nc22995, net_401}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc22996, nc22997, nc22998, nc22999, nc23000, nc23001, nc23002, nc23003, nc23004, nc23005, nc23006, nc23007, nc23008, nc23009, nc23010, nc23011, nc23012, nc23013, nc23014, nc23015, nc23016, nc23017, nc23018, nc23019, nc23020, nc23021, nc23022, nc23023, nc23024, nc23025, nc23026, nc23027, nc23028, nc23029, nc23030, nc23031, nc23032, nc23033, nc23034, nc23035, nc23036, nc23037, nc23038, nc23039, nc23040, nc23041, nc23042, nc23043, nc23044, nc23045, nc23046, nc23047, nc23048, nc23049, nc23050, nc23051, nc23052, nc23053, nc23054, nc23055, nc23056, nc23057, nc23058, dw[51]}),
		.dipa (),
		.dipb (),
		.cea (net_399),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_220 (
		.doa ({nc23059, nc23060, nc23061, nc23062, nc23063, nc23064, nc23065, nc23066, nc23067, nc23068, nc23069, nc23070, nc23071, nc23072, nc23073, nc23074, nc23075, nc23076, nc23077, nc23078, nc23079, nc23080, nc23081, nc23082, nc23083, nc23084, nc23085, nc23086, nc23087, nc23088, nc23089, nc23090, nc23091, nc23092, nc23093, nc23094, nc23095, nc23096, nc23097, nc23098, nc23099, nc23100, nc23101, nc23102, nc23103, nc23104, nc23105, nc23106, nc23107, nc23108, nc23109, nc23110, nc23111, nc23112, nc23113, nc23114, nc23115, nc23116, nc23117, nc23118, nc23119, nc23120, nc23121, net_405}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc23122, nc23123, nc23124, nc23125, nc23126, nc23127, nc23128, nc23129, nc23130, nc23131, nc23132, nc23133, nc23134, nc23135, nc23136, nc23137, nc23138, nc23139, nc23140, nc23141, nc23142, nc23143, nc23144, nc23145, nc23146, nc23147, nc23148, nc23149, nc23150, nc23151, nc23152, nc23153, nc23154, nc23155, nc23156, nc23157, nc23158, nc23159, nc23160, nc23161, nc23162, nc23163, nc23164, nc23165, nc23166, nc23167, nc23168, nc23169, nc23170, nc23171, nc23172, nc23173, nc23174, nc23175, nc23176, nc23177, nc23178, nc23179, nc23180, nc23181, nc23182, nc23183, nc23184, dw[59]}),
		.dipa (),
		.dipb (),
		.cea (net_403),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u196 (
		.sel (addra_pipe_0_net),
		.i0 (net_401),
		.i1 (net_405),
		.o (net_407)
	);
fifo2ram_emb_v1_AND u197 (
		.i0 (net_409),
		.i1 (net_408),
		.o (net_399)
	);
fifo2ram_emb_v1_AND u198 (
		.i0 (net_409),
		.i1 (ar[0]),
		.o (net_403)
	);
fifo2ram_emb_v1_NOT u199 (
		.i (ar[0]),
		.o (net_408)
	);
fifo2ram_emb_v1_MUX u200 (
		.sel (addra_pipe_1_net),
		.i0 (net_396),
		.i1 (net_407),
		.o (net_410)
	);
fifo2ram_emb_v1_AND u201 (
		.i0 (net_412),
		.i1 (net_411),
		.o (net_398)
	);
fifo2ram_emb_v1_AND u202 (
		.i0 (net_412),
		.i1 (ar[1]),
		.o (net_409)
	);
fifo2ram_emb_v1_NOT u203 (
		.i (ar[1]),
		.o (net_411)
	);
fifo2ram_emb_v1_MUX u204 (
		.sel (addra_pipe_2_net),
		.i0 (net_385),
		.i1 (net_410),
		.o (net_413)
	);
fifo2ram_emb_v1_AND u205 (
		.i0 (net_415),
		.i1 (net_414),
		.o (net_387)
	);
fifo2ram_emb_v1_AND u206 (
		.i0 (net_415),
		.i1 (ar[2]),
		.o (net_412)
	);
fifo2ram_emb_v1_NOT u207 (
		.i (ar[2]),
		.o (net_414)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_224 (
		.doa ({nc23185, nc23186, nc23187, nc23188, nc23189, nc23190, nc23191, nc23192, nc23193, nc23194, nc23195, nc23196, nc23197, nc23198, nc23199, nc23200, nc23201, nc23202, nc23203, nc23204, nc23205, nc23206, nc23207, nc23208, nc23209, nc23210, nc23211, nc23212, nc23213, nc23214, nc23215, nc23216, nc23217, nc23218, nc23219, nc23220, nc23221, nc23222, nc23223, nc23224, nc23225, nc23226, nc23227, nc23228, nc23229, nc23230, nc23231, nc23232, nc23233, nc23234, nc23235, nc23236, nc23237, nc23238, nc23239, nc23240, nc23241, nc23242, nc23243, nc23244, nc23245, nc23246, nc23247, net_418}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc23248, nc23249, nc23250, nc23251, nc23252, nc23253, nc23254, nc23255, nc23256, nc23257, nc23258, nc23259, nc23260, nc23261, nc23262, nc23263, nc23264, nc23265, nc23266, nc23267, nc23268, nc23269, nc23270, nc23271, nc23272, nc23273, nc23274, nc23275, nc23276, nc23277, nc23278, nc23279, nc23280, nc23281, nc23282, nc23283, nc23284, nc23285, nc23286, nc23287, nc23288, nc23289, nc23290, nc23291, nc23292, nc23293, nc23294, nc23295, nc23296, nc23297, nc23298, nc23299, nc23300, nc23301, nc23302, nc23303, nc23304, nc23305, nc23306, nc23307, nc23308, nc23309, nc23310, dw[67]}),
		.dipa (),
		.dipb (),
		.cea (net_416),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_228 (
		.doa ({nc23311, nc23312, nc23313, nc23314, nc23315, nc23316, nc23317, nc23318, nc23319, nc23320, nc23321, nc23322, nc23323, nc23324, nc23325, nc23326, nc23327, nc23328, nc23329, nc23330, nc23331, nc23332, nc23333, nc23334, nc23335, nc23336, nc23337, nc23338, nc23339, nc23340, nc23341, nc23342, nc23343, nc23344, nc23345, nc23346, nc23347, nc23348, nc23349, nc23350, nc23351, nc23352, nc23353, nc23354, nc23355, nc23356, nc23357, nc23358, nc23359, nc23360, nc23361, nc23362, nc23363, nc23364, nc23365, nc23366, nc23367, nc23368, nc23369, nc23370, nc23371, nc23372, nc23373, net_422}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc23374, nc23375, nc23376, nc23377, nc23378, nc23379, nc23380, nc23381, nc23382, nc23383, nc23384, nc23385, nc23386, nc23387, nc23388, nc23389, nc23390, nc23391, nc23392, nc23393, nc23394, nc23395, nc23396, nc23397, nc23398, nc23399, nc23400, nc23401, nc23402, nc23403, nc23404, nc23405, nc23406, nc23407, nc23408, nc23409, nc23410, nc23411, nc23412, nc23413, nc23414, nc23415, nc23416, nc23417, nc23418, nc23419, nc23420, nc23421, nc23422, nc23423, nc23424, nc23425, nc23426, nc23427, nc23428, nc23429, nc23430, nc23431, nc23432, nc23433, nc23434, nc23435, nc23436, dw[75]}),
		.dipa (),
		.dipb (),
		.cea (net_420),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u208 (
		.sel (addra_pipe_0_net),
		.i0 (net_418),
		.i1 (net_422),
		.o (net_424)
	);
fifo2ram_emb_v1_AND u209 (
		.i0 (net_426),
		.i1 (net_425),
		.o (net_416)
	);
fifo2ram_emb_v1_AND u210 (
		.i0 (net_426),
		.i1 (ar[0]),
		.o (net_420)
	);
fifo2ram_emb_v1_NOT u211 (
		.i (ar[0]),
		.o (net_425)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_232 (
		.doa ({nc23437, nc23438, nc23439, nc23440, nc23441, nc23442, nc23443, nc23444, nc23445, nc23446, nc23447, nc23448, nc23449, nc23450, nc23451, nc23452, nc23453, nc23454, nc23455, nc23456, nc23457, nc23458, nc23459, nc23460, nc23461, nc23462, nc23463, nc23464, nc23465, nc23466, nc23467, nc23468, nc23469, nc23470, nc23471, nc23472, nc23473, nc23474, nc23475, nc23476, nc23477, nc23478, nc23479, nc23480, nc23481, nc23482, nc23483, nc23484, nc23485, nc23486, nc23487, nc23488, nc23489, nc23490, nc23491, nc23492, nc23493, nc23494, nc23495, nc23496, nc23497, nc23498, nc23499, net_429}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc23500, nc23501, nc23502, nc23503, nc23504, nc23505, nc23506, nc23507, nc23508, nc23509, nc23510, nc23511, nc23512, nc23513, nc23514, nc23515, nc23516, nc23517, nc23518, nc23519, nc23520, nc23521, nc23522, nc23523, nc23524, nc23525, nc23526, nc23527, nc23528, nc23529, nc23530, nc23531, nc23532, nc23533, nc23534, nc23535, nc23536, nc23537, nc23538, nc23539, nc23540, nc23541, nc23542, nc23543, nc23544, nc23545, nc23546, nc23547, nc23548, nc23549, nc23550, nc23551, nc23552, nc23553, nc23554, nc23555, nc23556, nc23557, nc23558, nc23559, nc23560, nc23561, nc23562, dw[83]}),
		.dipa (),
		.dipb (),
		.cea (net_427),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_236 (
		.doa ({nc23563, nc23564, nc23565, nc23566, nc23567, nc23568, nc23569, nc23570, nc23571, nc23572, nc23573, nc23574, nc23575, nc23576, nc23577, nc23578, nc23579, nc23580, nc23581, nc23582, nc23583, nc23584, nc23585, nc23586, nc23587, nc23588, nc23589, nc23590, nc23591, nc23592, nc23593, nc23594, nc23595, nc23596, nc23597, nc23598, nc23599, nc23600, nc23601, nc23602, nc23603, nc23604, nc23605, nc23606, nc23607, nc23608, nc23609, nc23610, nc23611, nc23612, nc23613, nc23614, nc23615, nc23616, nc23617, nc23618, nc23619, nc23620, nc23621, nc23622, nc23623, nc23624, nc23625, net_433}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc23626, nc23627, nc23628, nc23629, nc23630, nc23631, nc23632, nc23633, nc23634, nc23635, nc23636, nc23637, nc23638, nc23639, nc23640, nc23641, nc23642, nc23643, nc23644, nc23645, nc23646, nc23647, nc23648, nc23649, nc23650, nc23651, nc23652, nc23653, nc23654, nc23655, nc23656, nc23657, nc23658, nc23659, nc23660, nc23661, nc23662, nc23663, nc23664, nc23665, nc23666, nc23667, nc23668, nc23669, nc23670, nc23671, nc23672, nc23673, nc23674, nc23675, nc23676, nc23677, nc23678, nc23679, nc23680, nc23681, nc23682, nc23683, nc23684, nc23685, nc23686, nc23687, nc23688, dw[91]}),
		.dipa (),
		.dipb (),
		.cea (net_431),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u212 (
		.sel (addra_pipe_0_net),
		.i0 (net_429),
		.i1 (net_433),
		.o (net_435)
	);
fifo2ram_emb_v1_AND u213 (
		.i0 (net_437),
		.i1 (net_436),
		.o (net_427)
	);
fifo2ram_emb_v1_AND u214 (
		.i0 (net_437),
		.i1 (ar[0]),
		.o (net_431)
	);
fifo2ram_emb_v1_NOT u215 (
		.i (ar[0]),
		.o (net_436)
	);
fifo2ram_emb_v1_MUX u216 (
		.sel (addra_pipe_1_net),
		.i0 (net_424),
		.i1 (net_435),
		.o (net_438)
	);
fifo2ram_emb_v1_AND u217 (
		.i0 (net_440),
		.i1 (net_439),
		.o (net_426)
	);
fifo2ram_emb_v1_AND u218 (
		.i0 (net_440),
		.i1 (ar[1]),
		.o (net_437)
	);
fifo2ram_emb_v1_NOT u219 (
		.i (ar[1]),
		.o (net_439)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_240 (
		.doa ({nc23689, nc23690, nc23691, nc23692, nc23693, nc23694, nc23695, nc23696, nc23697, nc23698, nc23699, nc23700, nc23701, nc23702, nc23703, nc23704, nc23705, nc23706, nc23707, nc23708, nc23709, nc23710, nc23711, nc23712, nc23713, nc23714, nc23715, nc23716, nc23717, nc23718, nc23719, nc23720, nc23721, nc23722, nc23723, nc23724, nc23725, nc23726, nc23727, nc23728, nc23729, nc23730, nc23731, nc23732, nc23733, nc23734, nc23735, nc23736, nc23737, nc23738, nc23739, nc23740, nc23741, nc23742, nc23743, nc23744, nc23745, nc23746, nc23747, nc23748, nc23749, nc23750, nc23751, net_443}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc23752, nc23753, nc23754, nc23755, nc23756, nc23757, nc23758, nc23759, nc23760, nc23761, nc23762, nc23763, nc23764, nc23765, nc23766, nc23767, nc23768, nc23769, nc23770, nc23771, nc23772, nc23773, nc23774, nc23775, nc23776, nc23777, nc23778, nc23779, nc23780, nc23781, nc23782, nc23783, nc23784, nc23785, nc23786, nc23787, nc23788, nc23789, nc23790, nc23791, nc23792, nc23793, nc23794, nc23795, nc23796, nc23797, nc23798, nc23799, nc23800, nc23801, nc23802, nc23803, nc23804, nc23805, nc23806, nc23807, nc23808, nc23809, nc23810, nc23811, nc23812, nc23813, nc23814, dw[99]}),
		.dipa (),
		.dipb (),
		.cea (net_441),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_244 (
		.doa ({nc23815, nc23816, nc23817, nc23818, nc23819, nc23820, nc23821, nc23822, nc23823, nc23824, nc23825, nc23826, nc23827, nc23828, nc23829, nc23830, nc23831, nc23832, nc23833, nc23834, nc23835, nc23836, nc23837, nc23838, nc23839, nc23840, nc23841, nc23842, nc23843, nc23844, nc23845, nc23846, nc23847, nc23848, nc23849, nc23850, nc23851, nc23852, nc23853, nc23854, nc23855, nc23856, nc23857, nc23858, nc23859, nc23860, nc23861, nc23862, nc23863, nc23864, nc23865, nc23866, nc23867, nc23868, nc23869, nc23870, nc23871, nc23872, nc23873, nc23874, nc23875, nc23876, nc23877, net_447}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc23878, nc23879, nc23880, nc23881, nc23882, nc23883, nc23884, nc23885, nc23886, nc23887, nc23888, nc23889, nc23890, nc23891, nc23892, nc23893, nc23894, nc23895, nc23896, nc23897, nc23898, nc23899, nc23900, nc23901, nc23902, nc23903, nc23904, nc23905, nc23906, nc23907, nc23908, nc23909, nc23910, nc23911, nc23912, nc23913, nc23914, nc23915, nc23916, nc23917, nc23918, nc23919, nc23920, nc23921, nc23922, nc23923, nc23924, nc23925, nc23926, nc23927, nc23928, nc23929, nc23930, nc23931, nc23932, nc23933, nc23934, nc23935, nc23936, nc23937, nc23938, nc23939, nc23940, dw[107]}),
		.dipa (),
		.dipb (),
		.cea (net_445),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u220 (
		.sel (addra_pipe_0_net),
		.i0 (net_443),
		.i1 (net_447),
		.o (net_449)
	);
fifo2ram_emb_v1_AND u221 (
		.i0 (net_451),
		.i1 (net_450),
		.o (net_441)
	);
fifo2ram_emb_v1_AND u222 (
		.i0 (net_451),
		.i1 (ar[0]),
		.o (net_445)
	);
fifo2ram_emb_v1_NOT u223 (
		.i (ar[0]),
		.o (net_450)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_248 (
		.doa ({nc23941, nc23942, nc23943, nc23944, nc23945, nc23946, nc23947, nc23948, nc23949, nc23950, nc23951, nc23952, nc23953, nc23954, nc23955, nc23956, nc23957, nc23958, nc23959, nc23960, nc23961, nc23962, nc23963, nc23964, nc23965, nc23966, nc23967, nc23968, nc23969, nc23970, nc23971, nc23972, nc23973, nc23974, nc23975, nc23976, nc23977, nc23978, nc23979, nc23980, nc23981, nc23982, nc23983, nc23984, nc23985, nc23986, nc23987, nc23988, nc23989, nc23990, nc23991, nc23992, nc23993, nc23994, nc23995, nc23996, nc23997, nc23998, nc23999, nc24000, nc24001, nc24002, nc24003, net_454}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24004, nc24005, nc24006, nc24007, nc24008, nc24009, nc24010, nc24011, nc24012, nc24013, nc24014, nc24015, nc24016, nc24017, nc24018, nc24019, nc24020, nc24021, nc24022, nc24023, nc24024, nc24025, nc24026, nc24027, nc24028, nc24029, nc24030, nc24031, nc24032, nc24033, nc24034, nc24035, nc24036, nc24037, nc24038, nc24039, nc24040, nc24041, nc24042, nc24043, nc24044, nc24045, nc24046, nc24047, nc24048, nc24049, nc24050, nc24051, nc24052, nc24053, nc24054, nc24055, nc24056, nc24057, nc24058, nc24059, nc24060, nc24061, nc24062, nc24063, nc24064, nc24065, nc24066, dw[115]}),
		.dipa (),
		.dipb (),
		.cea (net_452),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_252 (
		.doa ({nc24067, nc24068, nc24069, nc24070, nc24071, nc24072, nc24073, nc24074, nc24075, nc24076, nc24077, nc24078, nc24079, nc24080, nc24081, nc24082, nc24083, nc24084, nc24085, nc24086, nc24087, nc24088, nc24089, nc24090, nc24091, nc24092, nc24093, nc24094, nc24095, nc24096, nc24097, nc24098, nc24099, nc24100, nc24101, nc24102, nc24103, nc24104, nc24105, nc24106, nc24107, nc24108, nc24109, nc24110, nc24111, nc24112, nc24113, nc24114, nc24115, nc24116, nc24117, nc24118, nc24119, nc24120, nc24121, nc24122, nc24123, nc24124, nc24125, nc24126, nc24127, nc24128, nc24129, net_458}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24130, nc24131, nc24132, nc24133, nc24134, nc24135, nc24136, nc24137, nc24138, nc24139, nc24140, nc24141, nc24142, nc24143, nc24144, nc24145, nc24146, nc24147, nc24148, nc24149, nc24150, nc24151, nc24152, nc24153, nc24154, nc24155, nc24156, nc24157, nc24158, nc24159, nc24160, nc24161, nc24162, nc24163, nc24164, nc24165, nc24166, nc24167, nc24168, nc24169, nc24170, nc24171, nc24172, nc24173, nc24174, nc24175, nc24176, nc24177, nc24178, nc24179, nc24180, nc24181, nc24182, nc24183, nc24184, nc24185, nc24186, nc24187, nc24188, nc24189, nc24190, nc24191, nc24192, dw[123]}),
		.dipa (),
		.dipb (),
		.cea (net_456),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u224 (
		.sel (addra_pipe_0_net),
		.i0 (net_454),
		.i1 (net_458),
		.o (net_460)
	);
fifo2ram_emb_v1_AND u225 (
		.i0 (net_462),
		.i1 (net_461),
		.o (net_452)
	);
fifo2ram_emb_v1_AND u226 (
		.i0 (net_462),
		.i1 (ar[0]),
		.o (net_456)
	);
fifo2ram_emb_v1_NOT u227 (
		.i (ar[0]),
		.o (net_461)
	);
fifo2ram_emb_v1_MUX u228 (
		.sel (addra_pipe_1_net),
		.i0 (net_449),
		.i1 (net_460),
		.o (net_463)
	);
fifo2ram_emb_v1_AND u229 (
		.i0 (net_465),
		.i1 (net_464),
		.o (net_451)
	);
fifo2ram_emb_v1_AND u230 (
		.i0 (net_465),
		.i1 (ar[1]),
		.o (net_462)
	);
fifo2ram_emb_v1_NOT u231 (
		.i (ar[1]),
		.o (net_464)
	);
fifo2ram_emb_v1_MUX u232 (
		.sel (addra_pipe_2_net),
		.i0 (net_438),
		.i1 (net_463),
		.o (net_466)
	);
fifo2ram_emb_v1_AND u233 (
		.i0 (net_468),
		.i1 (net_467),
		.o (net_440)
	);
fifo2ram_emb_v1_AND u234 (
		.i0 (net_468),
		.i1 (ar[2]),
		.o (net_465)
	);
fifo2ram_emb_v1_NOT u235 (
		.i (ar[2]),
		.o (net_467)
	);
fifo2ram_emb_v1_MUX u236 (
		.sel (addra_pipe_3_net),
		.i0 (net_413),
		.i1 (net_466),
		.o (qr[3])
	);
fifo2ram_emb_v1_AND u237 (
		.i0 (cer),
		.i1 (net_470),
		.o (net_415)
	);
fifo2ram_emb_v1_AND u238 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_468)
	);
fifo2ram_emb_v1_NOT u239 (
		.i (ar[3]),
		.o (net_470)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_256 (
		.doa ({nc24193, nc24194, nc24195, nc24196, nc24197, nc24198, nc24199, nc24200, nc24201, nc24202, nc24203, nc24204, nc24205, nc24206, nc24207, nc24208, nc24209, nc24210, nc24211, nc24212, nc24213, nc24214, nc24215, nc24216, nc24217, nc24218, nc24219, nc24220, nc24221, nc24222, nc24223, nc24224, nc24225, nc24226, nc24227, nc24228, nc24229, nc24230, nc24231, nc24232, nc24233, nc24234, nc24235, nc24236, nc24237, nc24238, nc24239, nc24240, nc24241, nc24242, nc24243, nc24244, nc24245, nc24246, nc24247, nc24248, nc24249, nc24250, nc24251, nc24252, nc24253, nc24254, nc24255, net_474}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24256, nc24257, nc24258, nc24259, nc24260, nc24261, nc24262, nc24263, nc24264, nc24265, nc24266, nc24267, nc24268, nc24269, nc24270, nc24271, nc24272, nc24273, nc24274, nc24275, nc24276, nc24277, nc24278, nc24279, nc24280, nc24281, nc24282, nc24283, nc24284, nc24285, nc24286, nc24287, nc24288, nc24289, nc24290, nc24291, nc24292, nc24293, nc24294, nc24295, nc24296, nc24297, nc24298, nc24299, nc24300, nc24301, nc24302, nc24303, nc24304, nc24305, nc24306, nc24307, nc24308, nc24309, nc24310, nc24311, nc24312, nc24313, nc24314, nc24315, nc24316, nc24317, nc24318, dw[4]}),
		.dipa (),
		.dipb (),
		.cea (net_472),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_260 (
		.doa ({nc24319, nc24320, nc24321, nc24322, nc24323, nc24324, nc24325, nc24326, nc24327, nc24328, nc24329, nc24330, nc24331, nc24332, nc24333, nc24334, nc24335, nc24336, nc24337, nc24338, nc24339, nc24340, nc24341, nc24342, nc24343, nc24344, nc24345, nc24346, nc24347, nc24348, nc24349, nc24350, nc24351, nc24352, nc24353, nc24354, nc24355, nc24356, nc24357, nc24358, nc24359, nc24360, nc24361, nc24362, nc24363, nc24364, nc24365, nc24366, nc24367, nc24368, nc24369, nc24370, nc24371, nc24372, nc24373, nc24374, nc24375, nc24376, nc24377, nc24378, nc24379, nc24380, nc24381, net_478}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24382, nc24383, nc24384, nc24385, nc24386, nc24387, nc24388, nc24389, nc24390, nc24391, nc24392, nc24393, nc24394, nc24395, nc24396, nc24397, nc24398, nc24399, nc24400, nc24401, nc24402, nc24403, nc24404, nc24405, nc24406, nc24407, nc24408, nc24409, nc24410, nc24411, nc24412, nc24413, nc24414, nc24415, nc24416, nc24417, nc24418, nc24419, nc24420, nc24421, nc24422, nc24423, nc24424, nc24425, nc24426, nc24427, nc24428, nc24429, nc24430, nc24431, nc24432, nc24433, nc24434, nc24435, nc24436, nc24437, nc24438, nc24439, nc24440, nc24441, nc24442, nc24443, nc24444, dw[12]}),
		.dipa (),
		.dipb (),
		.cea (net_476),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u240 (
		.sel (addra_pipe_0_net),
		.i0 (net_474),
		.i1 (net_478),
		.o (net_480)
	);
fifo2ram_emb_v1_AND u241 (
		.i0 (net_482),
		.i1 (net_481),
		.o (net_472)
	);
fifo2ram_emb_v1_AND u242 (
		.i0 (net_482),
		.i1 (ar[0]),
		.o (net_476)
	);
fifo2ram_emb_v1_NOT u243 (
		.i (ar[0]),
		.o (net_481)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_264 (
		.doa ({nc24445, nc24446, nc24447, nc24448, nc24449, nc24450, nc24451, nc24452, nc24453, nc24454, nc24455, nc24456, nc24457, nc24458, nc24459, nc24460, nc24461, nc24462, nc24463, nc24464, nc24465, nc24466, nc24467, nc24468, nc24469, nc24470, nc24471, nc24472, nc24473, nc24474, nc24475, nc24476, nc24477, nc24478, nc24479, nc24480, nc24481, nc24482, nc24483, nc24484, nc24485, nc24486, nc24487, nc24488, nc24489, nc24490, nc24491, nc24492, nc24493, nc24494, nc24495, nc24496, nc24497, nc24498, nc24499, nc24500, nc24501, nc24502, nc24503, nc24504, nc24505, nc24506, nc24507, net_485}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24508, nc24509, nc24510, nc24511, nc24512, nc24513, nc24514, nc24515, nc24516, nc24517, nc24518, nc24519, nc24520, nc24521, nc24522, nc24523, nc24524, nc24525, nc24526, nc24527, nc24528, nc24529, nc24530, nc24531, nc24532, nc24533, nc24534, nc24535, nc24536, nc24537, nc24538, nc24539, nc24540, nc24541, nc24542, nc24543, nc24544, nc24545, nc24546, nc24547, nc24548, nc24549, nc24550, nc24551, nc24552, nc24553, nc24554, nc24555, nc24556, nc24557, nc24558, nc24559, nc24560, nc24561, nc24562, nc24563, nc24564, nc24565, nc24566, nc24567, nc24568, nc24569, nc24570, dw[20]}),
		.dipa (),
		.dipb (),
		.cea (net_483),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_268 (
		.doa ({nc24571, nc24572, nc24573, nc24574, nc24575, nc24576, nc24577, nc24578, nc24579, nc24580, nc24581, nc24582, nc24583, nc24584, nc24585, nc24586, nc24587, nc24588, nc24589, nc24590, nc24591, nc24592, nc24593, nc24594, nc24595, nc24596, nc24597, nc24598, nc24599, nc24600, nc24601, nc24602, nc24603, nc24604, nc24605, nc24606, nc24607, nc24608, nc24609, nc24610, nc24611, nc24612, nc24613, nc24614, nc24615, nc24616, nc24617, nc24618, nc24619, nc24620, nc24621, nc24622, nc24623, nc24624, nc24625, nc24626, nc24627, nc24628, nc24629, nc24630, nc24631, nc24632, nc24633, net_489}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24634, nc24635, nc24636, nc24637, nc24638, nc24639, nc24640, nc24641, nc24642, nc24643, nc24644, nc24645, nc24646, nc24647, nc24648, nc24649, nc24650, nc24651, nc24652, nc24653, nc24654, nc24655, nc24656, nc24657, nc24658, nc24659, nc24660, nc24661, nc24662, nc24663, nc24664, nc24665, nc24666, nc24667, nc24668, nc24669, nc24670, nc24671, nc24672, nc24673, nc24674, nc24675, nc24676, nc24677, nc24678, nc24679, nc24680, nc24681, nc24682, nc24683, nc24684, nc24685, nc24686, nc24687, nc24688, nc24689, nc24690, nc24691, nc24692, nc24693, nc24694, nc24695, nc24696, dw[28]}),
		.dipa (),
		.dipb (),
		.cea (net_487),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u244 (
		.sel (addra_pipe_0_net),
		.i0 (net_485),
		.i1 (net_489),
		.o (net_491)
	);
fifo2ram_emb_v1_AND u245 (
		.i0 (net_493),
		.i1 (net_492),
		.o (net_483)
	);
fifo2ram_emb_v1_AND u246 (
		.i0 (net_493),
		.i1 (ar[0]),
		.o (net_487)
	);
fifo2ram_emb_v1_NOT u247 (
		.i (ar[0]),
		.o (net_492)
	);
fifo2ram_emb_v1_MUX u248 (
		.sel (addra_pipe_1_net),
		.i0 (net_480),
		.i1 (net_491),
		.o (net_494)
	);
fifo2ram_emb_v1_AND u249 (
		.i0 (net_496),
		.i1 (net_495),
		.o (net_482)
	);
fifo2ram_emb_v1_AND u250 (
		.i0 (net_496),
		.i1 (ar[1]),
		.o (net_493)
	);
fifo2ram_emb_v1_NOT u251 (
		.i (ar[1]),
		.o (net_495)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_272 (
		.doa ({nc24697, nc24698, nc24699, nc24700, nc24701, nc24702, nc24703, nc24704, nc24705, nc24706, nc24707, nc24708, nc24709, nc24710, nc24711, nc24712, nc24713, nc24714, nc24715, nc24716, nc24717, nc24718, nc24719, nc24720, nc24721, nc24722, nc24723, nc24724, nc24725, nc24726, nc24727, nc24728, nc24729, nc24730, nc24731, nc24732, nc24733, nc24734, nc24735, nc24736, nc24737, nc24738, nc24739, nc24740, nc24741, nc24742, nc24743, nc24744, nc24745, nc24746, nc24747, nc24748, nc24749, nc24750, nc24751, nc24752, nc24753, nc24754, nc24755, nc24756, nc24757, nc24758, nc24759, net_499}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24760, nc24761, nc24762, nc24763, nc24764, nc24765, nc24766, nc24767, nc24768, nc24769, nc24770, nc24771, nc24772, nc24773, nc24774, nc24775, nc24776, nc24777, nc24778, nc24779, nc24780, nc24781, nc24782, nc24783, nc24784, nc24785, nc24786, nc24787, nc24788, nc24789, nc24790, nc24791, nc24792, nc24793, nc24794, nc24795, nc24796, nc24797, nc24798, nc24799, nc24800, nc24801, nc24802, nc24803, nc24804, nc24805, nc24806, nc24807, nc24808, nc24809, nc24810, nc24811, nc24812, nc24813, nc24814, nc24815, nc24816, nc24817, nc24818, nc24819, nc24820, nc24821, nc24822, dw[36]}),
		.dipa (),
		.dipb (),
		.cea (net_497),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_276 (
		.doa ({nc24823, nc24824, nc24825, nc24826, nc24827, nc24828, nc24829, nc24830, nc24831, nc24832, nc24833, nc24834, nc24835, nc24836, nc24837, nc24838, nc24839, nc24840, nc24841, nc24842, nc24843, nc24844, nc24845, nc24846, nc24847, nc24848, nc24849, nc24850, nc24851, nc24852, nc24853, nc24854, nc24855, nc24856, nc24857, nc24858, nc24859, nc24860, nc24861, nc24862, nc24863, nc24864, nc24865, nc24866, nc24867, nc24868, nc24869, nc24870, nc24871, nc24872, nc24873, nc24874, nc24875, nc24876, nc24877, nc24878, nc24879, nc24880, nc24881, nc24882, nc24883, nc24884, nc24885, net_503}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc24886, nc24887, nc24888, nc24889, nc24890, nc24891, nc24892, nc24893, nc24894, nc24895, nc24896, nc24897, nc24898, nc24899, nc24900, nc24901, nc24902, nc24903, nc24904, nc24905, nc24906, nc24907, nc24908, nc24909, nc24910, nc24911, nc24912, nc24913, nc24914, nc24915, nc24916, nc24917, nc24918, nc24919, nc24920, nc24921, nc24922, nc24923, nc24924, nc24925, nc24926, nc24927, nc24928, nc24929, nc24930, nc24931, nc24932, nc24933, nc24934, nc24935, nc24936, nc24937, nc24938, nc24939, nc24940, nc24941, nc24942, nc24943, nc24944, nc24945, nc24946, nc24947, nc24948, dw[44]}),
		.dipa (),
		.dipb (),
		.cea (net_501),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u252 (
		.sel (addra_pipe_0_net),
		.i0 (net_499),
		.i1 (net_503),
		.o (net_505)
	);
fifo2ram_emb_v1_AND u253 (
		.i0 (net_507),
		.i1 (net_506),
		.o (net_497)
	);
fifo2ram_emb_v1_AND u254 (
		.i0 (net_507),
		.i1 (ar[0]),
		.o (net_501)
	);
fifo2ram_emb_v1_NOT u255 (
		.i (ar[0]),
		.o (net_506)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_280 (
		.doa ({nc24949, nc24950, nc24951, nc24952, nc24953, nc24954, nc24955, nc24956, nc24957, nc24958, nc24959, nc24960, nc24961, nc24962, nc24963, nc24964, nc24965, nc24966, nc24967, nc24968, nc24969, nc24970, nc24971, nc24972, nc24973, nc24974, nc24975, nc24976, nc24977, nc24978, nc24979, nc24980, nc24981, nc24982, nc24983, nc24984, nc24985, nc24986, nc24987, nc24988, nc24989, nc24990, nc24991, nc24992, nc24993, nc24994, nc24995, nc24996, nc24997, nc24998, nc24999, nc25000, nc25001, nc25002, nc25003, nc25004, nc25005, nc25006, nc25007, nc25008, nc25009, nc25010, nc25011, net_510}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25012, nc25013, nc25014, nc25015, nc25016, nc25017, nc25018, nc25019, nc25020, nc25021, nc25022, nc25023, nc25024, nc25025, nc25026, nc25027, nc25028, nc25029, nc25030, nc25031, nc25032, nc25033, nc25034, nc25035, nc25036, nc25037, nc25038, nc25039, nc25040, nc25041, nc25042, nc25043, nc25044, nc25045, nc25046, nc25047, nc25048, nc25049, nc25050, nc25051, nc25052, nc25053, nc25054, nc25055, nc25056, nc25057, nc25058, nc25059, nc25060, nc25061, nc25062, nc25063, nc25064, nc25065, nc25066, nc25067, nc25068, nc25069, nc25070, nc25071, nc25072, nc25073, nc25074, dw[52]}),
		.dipa (),
		.dipb (),
		.cea (net_508),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_284 (
		.doa ({nc25075, nc25076, nc25077, nc25078, nc25079, nc25080, nc25081, nc25082, nc25083, nc25084, nc25085, nc25086, nc25087, nc25088, nc25089, nc25090, nc25091, nc25092, nc25093, nc25094, nc25095, nc25096, nc25097, nc25098, nc25099, nc25100, nc25101, nc25102, nc25103, nc25104, nc25105, nc25106, nc25107, nc25108, nc25109, nc25110, nc25111, nc25112, nc25113, nc25114, nc25115, nc25116, nc25117, nc25118, nc25119, nc25120, nc25121, nc25122, nc25123, nc25124, nc25125, nc25126, nc25127, nc25128, nc25129, nc25130, nc25131, nc25132, nc25133, nc25134, nc25135, nc25136, nc25137, net_514}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25138, nc25139, nc25140, nc25141, nc25142, nc25143, nc25144, nc25145, nc25146, nc25147, nc25148, nc25149, nc25150, nc25151, nc25152, nc25153, nc25154, nc25155, nc25156, nc25157, nc25158, nc25159, nc25160, nc25161, nc25162, nc25163, nc25164, nc25165, nc25166, nc25167, nc25168, nc25169, nc25170, nc25171, nc25172, nc25173, nc25174, nc25175, nc25176, nc25177, nc25178, nc25179, nc25180, nc25181, nc25182, nc25183, nc25184, nc25185, nc25186, nc25187, nc25188, nc25189, nc25190, nc25191, nc25192, nc25193, nc25194, nc25195, nc25196, nc25197, nc25198, nc25199, nc25200, dw[60]}),
		.dipa (),
		.dipb (),
		.cea (net_512),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u256 (
		.sel (addra_pipe_0_net),
		.i0 (net_510),
		.i1 (net_514),
		.o (net_516)
	);
fifo2ram_emb_v1_AND u257 (
		.i0 (net_518),
		.i1 (net_517),
		.o (net_508)
	);
fifo2ram_emb_v1_AND u258 (
		.i0 (net_518),
		.i1 (ar[0]),
		.o (net_512)
	);
fifo2ram_emb_v1_NOT u259 (
		.i (ar[0]),
		.o (net_517)
	);
fifo2ram_emb_v1_MUX u260 (
		.sel (addra_pipe_1_net),
		.i0 (net_505),
		.i1 (net_516),
		.o (net_519)
	);
fifo2ram_emb_v1_AND u261 (
		.i0 (net_521),
		.i1 (net_520),
		.o (net_507)
	);
fifo2ram_emb_v1_AND u262 (
		.i0 (net_521),
		.i1 (ar[1]),
		.o (net_518)
	);
fifo2ram_emb_v1_NOT u263 (
		.i (ar[1]),
		.o (net_520)
	);
fifo2ram_emb_v1_MUX u264 (
		.sel (addra_pipe_2_net),
		.i0 (net_494),
		.i1 (net_519),
		.o (net_522)
	);
fifo2ram_emb_v1_AND u265 (
		.i0 (net_524),
		.i1 (net_523),
		.o (net_496)
	);
fifo2ram_emb_v1_AND u266 (
		.i0 (net_524),
		.i1 (ar[2]),
		.o (net_521)
	);
fifo2ram_emb_v1_NOT u267 (
		.i (ar[2]),
		.o (net_523)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_288 (
		.doa ({nc25201, nc25202, nc25203, nc25204, nc25205, nc25206, nc25207, nc25208, nc25209, nc25210, nc25211, nc25212, nc25213, nc25214, nc25215, nc25216, nc25217, nc25218, nc25219, nc25220, nc25221, nc25222, nc25223, nc25224, nc25225, nc25226, nc25227, nc25228, nc25229, nc25230, nc25231, nc25232, nc25233, nc25234, nc25235, nc25236, nc25237, nc25238, nc25239, nc25240, nc25241, nc25242, nc25243, nc25244, nc25245, nc25246, nc25247, nc25248, nc25249, nc25250, nc25251, nc25252, nc25253, nc25254, nc25255, nc25256, nc25257, nc25258, nc25259, nc25260, nc25261, nc25262, nc25263, net_527}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25264, nc25265, nc25266, nc25267, nc25268, nc25269, nc25270, nc25271, nc25272, nc25273, nc25274, nc25275, nc25276, nc25277, nc25278, nc25279, nc25280, nc25281, nc25282, nc25283, nc25284, nc25285, nc25286, nc25287, nc25288, nc25289, nc25290, nc25291, nc25292, nc25293, nc25294, nc25295, nc25296, nc25297, nc25298, nc25299, nc25300, nc25301, nc25302, nc25303, nc25304, nc25305, nc25306, nc25307, nc25308, nc25309, nc25310, nc25311, nc25312, nc25313, nc25314, nc25315, nc25316, nc25317, nc25318, nc25319, nc25320, nc25321, nc25322, nc25323, nc25324, nc25325, nc25326, dw[68]}),
		.dipa (),
		.dipb (),
		.cea (net_525),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_292 (
		.doa ({nc25327, nc25328, nc25329, nc25330, nc25331, nc25332, nc25333, nc25334, nc25335, nc25336, nc25337, nc25338, nc25339, nc25340, nc25341, nc25342, nc25343, nc25344, nc25345, nc25346, nc25347, nc25348, nc25349, nc25350, nc25351, nc25352, nc25353, nc25354, nc25355, nc25356, nc25357, nc25358, nc25359, nc25360, nc25361, nc25362, nc25363, nc25364, nc25365, nc25366, nc25367, nc25368, nc25369, nc25370, nc25371, nc25372, nc25373, nc25374, nc25375, nc25376, nc25377, nc25378, nc25379, nc25380, nc25381, nc25382, nc25383, nc25384, nc25385, nc25386, nc25387, nc25388, nc25389, net_531}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25390, nc25391, nc25392, nc25393, nc25394, nc25395, nc25396, nc25397, nc25398, nc25399, nc25400, nc25401, nc25402, nc25403, nc25404, nc25405, nc25406, nc25407, nc25408, nc25409, nc25410, nc25411, nc25412, nc25413, nc25414, nc25415, nc25416, nc25417, nc25418, nc25419, nc25420, nc25421, nc25422, nc25423, nc25424, nc25425, nc25426, nc25427, nc25428, nc25429, nc25430, nc25431, nc25432, nc25433, nc25434, nc25435, nc25436, nc25437, nc25438, nc25439, nc25440, nc25441, nc25442, nc25443, nc25444, nc25445, nc25446, nc25447, nc25448, nc25449, nc25450, nc25451, nc25452, dw[76]}),
		.dipa (),
		.dipb (),
		.cea (net_529),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u268 (
		.sel (addra_pipe_0_net),
		.i0 (net_527),
		.i1 (net_531),
		.o (net_533)
	);
fifo2ram_emb_v1_AND u269 (
		.i0 (net_535),
		.i1 (net_534),
		.o (net_525)
	);
fifo2ram_emb_v1_AND u270 (
		.i0 (net_535),
		.i1 (ar[0]),
		.o (net_529)
	);
fifo2ram_emb_v1_NOT u271 (
		.i (ar[0]),
		.o (net_534)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_296 (
		.doa ({nc25453, nc25454, nc25455, nc25456, nc25457, nc25458, nc25459, nc25460, nc25461, nc25462, nc25463, nc25464, nc25465, nc25466, nc25467, nc25468, nc25469, nc25470, nc25471, nc25472, nc25473, nc25474, nc25475, nc25476, nc25477, nc25478, nc25479, nc25480, nc25481, nc25482, nc25483, nc25484, nc25485, nc25486, nc25487, nc25488, nc25489, nc25490, nc25491, nc25492, nc25493, nc25494, nc25495, nc25496, nc25497, nc25498, nc25499, nc25500, nc25501, nc25502, nc25503, nc25504, nc25505, nc25506, nc25507, nc25508, nc25509, nc25510, nc25511, nc25512, nc25513, nc25514, nc25515, net_538}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25516, nc25517, nc25518, nc25519, nc25520, nc25521, nc25522, nc25523, nc25524, nc25525, nc25526, nc25527, nc25528, nc25529, nc25530, nc25531, nc25532, nc25533, nc25534, nc25535, nc25536, nc25537, nc25538, nc25539, nc25540, nc25541, nc25542, nc25543, nc25544, nc25545, nc25546, nc25547, nc25548, nc25549, nc25550, nc25551, nc25552, nc25553, nc25554, nc25555, nc25556, nc25557, nc25558, nc25559, nc25560, nc25561, nc25562, nc25563, nc25564, nc25565, nc25566, nc25567, nc25568, nc25569, nc25570, nc25571, nc25572, nc25573, nc25574, nc25575, nc25576, nc25577, nc25578, dw[84]}),
		.dipa (),
		.dipb (),
		.cea (net_536),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_300 (
		.doa ({nc25579, nc25580, nc25581, nc25582, nc25583, nc25584, nc25585, nc25586, nc25587, nc25588, nc25589, nc25590, nc25591, nc25592, nc25593, nc25594, nc25595, nc25596, nc25597, nc25598, nc25599, nc25600, nc25601, nc25602, nc25603, nc25604, nc25605, nc25606, nc25607, nc25608, nc25609, nc25610, nc25611, nc25612, nc25613, nc25614, nc25615, nc25616, nc25617, nc25618, nc25619, nc25620, nc25621, nc25622, nc25623, nc25624, nc25625, nc25626, nc25627, nc25628, nc25629, nc25630, nc25631, nc25632, nc25633, nc25634, nc25635, nc25636, nc25637, nc25638, nc25639, nc25640, nc25641, net_542}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25642, nc25643, nc25644, nc25645, nc25646, nc25647, nc25648, nc25649, nc25650, nc25651, nc25652, nc25653, nc25654, nc25655, nc25656, nc25657, nc25658, nc25659, nc25660, nc25661, nc25662, nc25663, nc25664, nc25665, nc25666, nc25667, nc25668, nc25669, nc25670, nc25671, nc25672, nc25673, nc25674, nc25675, nc25676, nc25677, nc25678, nc25679, nc25680, nc25681, nc25682, nc25683, nc25684, nc25685, nc25686, nc25687, nc25688, nc25689, nc25690, nc25691, nc25692, nc25693, nc25694, nc25695, nc25696, nc25697, nc25698, nc25699, nc25700, nc25701, nc25702, nc25703, nc25704, dw[92]}),
		.dipa (),
		.dipb (),
		.cea (net_540),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u272 (
		.sel (addra_pipe_0_net),
		.i0 (net_538),
		.i1 (net_542),
		.o (net_544)
	);
fifo2ram_emb_v1_AND u273 (
		.i0 (net_546),
		.i1 (net_545),
		.o (net_536)
	);
fifo2ram_emb_v1_AND u274 (
		.i0 (net_546),
		.i1 (ar[0]),
		.o (net_540)
	);
fifo2ram_emb_v1_NOT u275 (
		.i (ar[0]),
		.o (net_545)
	);
fifo2ram_emb_v1_MUX u276 (
		.sel (addra_pipe_1_net),
		.i0 (net_533),
		.i1 (net_544),
		.o (net_547)
	);
fifo2ram_emb_v1_AND u277 (
		.i0 (net_549),
		.i1 (net_548),
		.o (net_535)
	);
fifo2ram_emb_v1_AND u278 (
		.i0 (net_549),
		.i1 (ar[1]),
		.o (net_546)
	);
fifo2ram_emb_v1_NOT u279 (
		.i (ar[1]),
		.o (net_548)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_304 (
		.doa ({nc25705, nc25706, nc25707, nc25708, nc25709, nc25710, nc25711, nc25712, nc25713, nc25714, nc25715, nc25716, nc25717, nc25718, nc25719, nc25720, nc25721, nc25722, nc25723, nc25724, nc25725, nc25726, nc25727, nc25728, nc25729, nc25730, nc25731, nc25732, nc25733, nc25734, nc25735, nc25736, nc25737, nc25738, nc25739, nc25740, nc25741, nc25742, nc25743, nc25744, nc25745, nc25746, nc25747, nc25748, nc25749, nc25750, nc25751, nc25752, nc25753, nc25754, nc25755, nc25756, nc25757, nc25758, nc25759, nc25760, nc25761, nc25762, nc25763, nc25764, nc25765, nc25766, nc25767, net_552}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25768, nc25769, nc25770, nc25771, nc25772, nc25773, nc25774, nc25775, nc25776, nc25777, nc25778, nc25779, nc25780, nc25781, nc25782, nc25783, nc25784, nc25785, nc25786, nc25787, nc25788, nc25789, nc25790, nc25791, nc25792, nc25793, nc25794, nc25795, nc25796, nc25797, nc25798, nc25799, nc25800, nc25801, nc25802, nc25803, nc25804, nc25805, nc25806, nc25807, nc25808, nc25809, nc25810, nc25811, nc25812, nc25813, nc25814, nc25815, nc25816, nc25817, nc25818, nc25819, nc25820, nc25821, nc25822, nc25823, nc25824, nc25825, nc25826, nc25827, nc25828, nc25829, nc25830, dw[100]}),
		.dipa (),
		.dipb (),
		.cea (net_550),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_308 (
		.doa ({nc25831, nc25832, nc25833, nc25834, nc25835, nc25836, nc25837, nc25838, nc25839, nc25840, nc25841, nc25842, nc25843, nc25844, nc25845, nc25846, nc25847, nc25848, nc25849, nc25850, nc25851, nc25852, nc25853, nc25854, nc25855, nc25856, nc25857, nc25858, nc25859, nc25860, nc25861, nc25862, nc25863, nc25864, nc25865, nc25866, nc25867, nc25868, nc25869, nc25870, nc25871, nc25872, nc25873, nc25874, nc25875, nc25876, nc25877, nc25878, nc25879, nc25880, nc25881, nc25882, nc25883, nc25884, nc25885, nc25886, nc25887, nc25888, nc25889, nc25890, nc25891, nc25892, nc25893, net_556}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc25894, nc25895, nc25896, nc25897, nc25898, nc25899, nc25900, nc25901, nc25902, nc25903, nc25904, nc25905, nc25906, nc25907, nc25908, nc25909, nc25910, nc25911, nc25912, nc25913, nc25914, nc25915, nc25916, nc25917, nc25918, nc25919, nc25920, nc25921, nc25922, nc25923, nc25924, nc25925, nc25926, nc25927, nc25928, nc25929, nc25930, nc25931, nc25932, nc25933, nc25934, nc25935, nc25936, nc25937, nc25938, nc25939, nc25940, nc25941, nc25942, nc25943, nc25944, nc25945, nc25946, nc25947, nc25948, nc25949, nc25950, nc25951, nc25952, nc25953, nc25954, nc25955, nc25956, dw[108]}),
		.dipa (),
		.dipb (),
		.cea (net_554),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u280 (
		.sel (addra_pipe_0_net),
		.i0 (net_552),
		.i1 (net_556),
		.o (net_558)
	);
fifo2ram_emb_v1_AND u281 (
		.i0 (net_560),
		.i1 (net_559),
		.o (net_550)
	);
fifo2ram_emb_v1_AND u282 (
		.i0 (net_560),
		.i1 (ar[0]),
		.o (net_554)
	);
fifo2ram_emb_v1_NOT u283 (
		.i (ar[0]),
		.o (net_559)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_312 (
		.doa ({nc25957, nc25958, nc25959, nc25960, nc25961, nc25962, nc25963, nc25964, nc25965, nc25966, nc25967, nc25968, nc25969, nc25970, nc25971, nc25972, nc25973, nc25974, nc25975, nc25976, nc25977, nc25978, nc25979, nc25980, nc25981, nc25982, nc25983, nc25984, nc25985, nc25986, nc25987, nc25988, nc25989, nc25990, nc25991, nc25992, nc25993, nc25994, nc25995, nc25996, nc25997, nc25998, nc25999, nc26000, nc26001, nc26002, nc26003, nc26004, nc26005, nc26006, nc26007, nc26008, nc26009, nc26010, nc26011, nc26012, nc26013, nc26014, nc26015, nc26016, nc26017, nc26018, nc26019, net_563}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26020, nc26021, nc26022, nc26023, nc26024, nc26025, nc26026, nc26027, nc26028, nc26029, nc26030, nc26031, nc26032, nc26033, nc26034, nc26035, nc26036, nc26037, nc26038, nc26039, nc26040, nc26041, nc26042, nc26043, nc26044, nc26045, nc26046, nc26047, nc26048, nc26049, nc26050, nc26051, nc26052, nc26053, nc26054, nc26055, nc26056, nc26057, nc26058, nc26059, nc26060, nc26061, nc26062, nc26063, nc26064, nc26065, nc26066, nc26067, nc26068, nc26069, nc26070, nc26071, nc26072, nc26073, nc26074, nc26075, nc26076, nc26077, nc26078, nc26079, nc26080, nc26081, nc26082, dw[116]}),
		.dipa (),
		.dipb (),
		.cea (net_561),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_316 (
		.doa ({nc26083, nc26084, nc26085, nc26086, nc26087, nc26088, nc26089, nc26090, nc26091, nc26092, nc26093, nc26094, nc26095, nc26096, nc26097, nc26098, nc26099, nc26100, nc26101, nc26102, nc26103, nc26104, nc26105, nc26106, nc26107, nc26108, nc26109, nc26110, nc26111, nc26112, nc26113, nc26114, nc26115, nc26116, nc26117, nc26118, nc26119, nc26120, nc26121, nc26122, nc26123, nc26124, nc26125, nc26126, nc26127, nc26128, nc26129, nc26130, nc26131, nc26132, nc26133, nc26134, nc26135, nc26136, nc26137, nc26138, nc26139, nc26140, nc26141, nc26142, nc26143, nc26144, nc26145, net_567}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26146, nc26147, nc26148, nc26149, nc26150, nc26151, nc26152, nc26153, nc26154, nc26155, nc26156, nc26157, nc26158, nc26159, nc26160, nc26161, nc26162, nc26163, nc26164, nc26165, nc26166, nc26167, nc26168, nc26169, nc26170, nc26171, nc26172, nc26173, nc26174, nc26175, nc26176, nc26177, nc26178, nc26179, nc26180, nc26181, nc26182, nc26183, nc26184, nc26185, nc26186, nc26187, nc26188, nc26189, nc26190, nc26191, nc26192, nc26193, nc26194, nc26195, nc26196, nc26197, nc26198, nc26199, nc26200, nc26201, nc26202, nc26203, nc26204, nc26205, nc26206, nc26207, nc26208, dw[124]}),
		.dipa (),
		.dipb (),
		.cea (net_565),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u284 (
		.sel (addra_pipe_0_net),
		.i0 (net_563),
		.i1 (net_567),
		.o (net_569)
	);
fifo2ram_emb_v1_AND u285 (
		.i0 (net_571),
		.i1 (net_570),
		.o (net_561)
	);
fifo2ram_emb_v1_AND u286 (
		.i0 (net_571),
		.i1 (ar[0]),
		.o (net_565)
	);
fifo2ram_emb_v1_NOT u287 (
		.i (ar[0]),
		.o (net_570)
	);
fifo2ram_emb_v1_MUX u288 (
		.sel (addra_pipe_1_net),
		.i0 (net_558),
		.i1 (net_569),
		.o (net_572)
	);
fifo2ram_emb_v1_AND u289 (
		.i0 (net_574),
		.i1 (net_573),
		.o (net_560)
	);
fifo2ram_emb_v1_AND u290 (
		.i0 (net_574),
		.i1 (ar[1]),
		.o (net_571)
	);
fifo2ram_emb_v1_NOT u291 (
		.i (ar[1]),
		.o (net_573)
	);
fifo2ram_emb_v1_MUX u292 (
		.sel (addra_pipe_2_net),
		.i0 (net_547),
		.i1 (net_572),
		.o (net_575)
	);
fifo2ram_emb_v1_AND u293 (
		.i0 (net_577),
		.i1 (net_576),
		.o (net_549)
	);
fifo2ram_emb_v1_AND u294 (
		.i0 (net_577),
		.i1 (ar[2]),
		.o (net_574)
	);
fifo2ram_emb_v1_NOT u295 (
		.i (ar[2]),
		.o (net_576)
	);
fifo2ram_emb_v1_MUX u296 (
		.sel (addra_pipe_3_net),
		.i0 (net_522),
		.i1 (net_575),
		.o (qr[4])
	);
fifo2ram_emb_v1_AND u297 (
		.i0 (cer),
		.i1 (net_579),
		.o (net_524)
	);
fifo2ram_emb_v1_AND u298 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_577)
	);
fifo2ram_emb_v1_NOT u299 (
		.i (ar[3]),
		.o (net_579)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_320 (
		.doa ({nc26209, nc26210, nc26211, nc26212, nc26213, nc26214, nc26215, nc26216, nc26217, nc26218, nc26219, nc26220, nc26221, nc26222, nc26223, nc26224, nc26225, nc26226, nc26227, nc26228, nc26229, nc26230, nc26231, nc26232, nc26233, nc26234, nc26235, nc26236, nc26237, nc26238, nc26239, nc26240, nc26241, nc26242, nc26243, nc26244, nc26245, nc26246, nc26247, nc26248, nc26249, nc26250, nc26251, nc26252, nc26253, nc26254, nc26255, nc26256, nc26257, nc26258, nc26259, nc26260, nc26261, nc26262, nc26263, nc26264, nc26265, nc26266, nc26267, nc26268, nc26269, nc26270, nc26271, net_583}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26272, nc26273, nc26274, nc26275, nc26276, nc26277, nc26278, nc26279, nc26280, nc26281, nc26282, nc26283, nc26284, nc26285, nc26286, nc26287, nc26288, nc26289, nc26290, nc26291, nc26292, nc26293, nc26294, nc26295, nc26296, nc26297, nc26298, nc26299, nc26300, nc26301, nc26302, nc26303, nc26304, nc26305, nc26306, nc26307, nc26308, nc26309, nc26310, nc26311, nc26312, nc26313, nc26314, nc26315, nc26316, nc26317, nc26318, nc26319, nc26320, nc26321, nc26322, nc26323, nc26324, nc26325, nc26326, nc26327, nc26328, nc26329, nc26330, nc26331, nc26332, nc26333, nc26334, dw[5]}),
		.dipa (),
		.dipb (),
		.cea (net_581),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_324 (
		.doa ({nc26335, nc26336, nc26337, nc26338, nc26339, nc26340, nc26341, nc26342, nc26343, nc26344, nc26345, nc26346, nc26347, nc26348, nc26349, nc26350, nc26351, nc26352, nc26353, nc26354, nc26355, nc26356, nc26357, nc26358, nc26359, nc26360, nc26361, nc26362, nc26363, nc26364, nc26365, nc26366, nc26367, nc26368, nc26369, nc26370, nc26371, nc26372, nc26373, nc26374, nc26375, nc26376, nc26377, nc26378, nc26379, nc26380, nc26381, nc26382, nc26383, nc26384, nc26385, nc26386, nc26387, nc26388, nc26389, nc26390, nc26391, nc26392, nc26393, nc26394, nc26395, nc26396, nc26397, net_587}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26398, nc26399, nc26400, nc26401, nc26402, nc26403, nc26404, nc26405, nc26406, nc26407, nc26408, nc26409, nc26410, nc26411, nc26412, nc26413, nc26414, nc26415, nc26416, nc26417, nc26418, nc26419, nc26420, nc26421, nc26422, nc26423, nc26424, nc26425, nc26426, nc26427, nc26428, nc26429, nc26430, nc26431, nc26432, nc26433, nc26434, nc26435, nc26436, nc26437, nc26438, nc26439, nc26440, nc26441, nc26442, nc26443, nc26444, nc26445, nc26446, nc26447, nc26448, nc26449, nc26450, nc26451, nc26452, nc26453, nc26454, nc26455, nc26456, nc26457, nc26458, nc26459, nc26460, dw[13]}),
		.dipa (),
		.dipb (),
		.cea (net_585),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u300 (
		.sel (addra_pipe_0_net),
		.i0 (net_583),
		.i1 (net_587),
		.o (net_589)
	);
fifo2ram_emb_v1_AND u301 (
		.i0 (net_591),
		.i1 (net_590),
		.o (net_581)
	);
fifo2ram_emb_v1_AND u302 (
		.i0 (net_591),
		.i1 (ar[0]),
		.o (net_585)
	);
fifo2ram_emb_v1_NOT u303 (
		.i (ar[0]),
		.o (net_590)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_328 (
		.doa ({nc26461, nc26462, nc26463, nc26464, nc26465, nc26466, nc26467, nc26468, nc26469, nc26470, nc26471, nc26472, nc26473, nc26474, nc26475, nc26476, nc26477, nc26478, nc26479, nc26480, nc26481, nc26482, nc26483, nc26484, nc26485, nc26486, nc26487, nc26488, nc26489, nc26490, nc26491, nc26492, nc26493, nc26494, nc26495, nc26496, nc26497, nc26498, nc26499, nc26500, nc26501, nc26502, nc26503, nc26504, nc26505, nc26506, nc26507, nc26508, nc26509, nc26510, nc26511, nc26512, nc26513, nc26514, nc26515, nc26516, nc26517, nc26518, nc26519, nc26520, nc26521, nc26522, nc26523, net_594}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26524, nc26525, nc26526, nc26527, nc26528, nc26529, nc26530, nc26531, nc26532, nc26533, nc26534, nc26535, nc26536, nc26537, nc26538, nc26539, nc26540, nc26541, nc26542, nc26543, nc26544, nc26545, nc26546, nc26547, nc26548, nc26549, nc26550, nc26551, nc26552, nc26553, nc26554, nc26555, nc26556, nc26557, nc26558, nc26559, nc26560, nc26561, nc26562, nc26563, nc26564, nc26565, nc26566, nc26567, nc26568, nc26569, nc26570, nc26571, nc26572, nc26573, nc26574, nc26575, nc26576, nc26577, nc26578, nc26579, nc26580, nc26581, nc26582, nc26583, nc26584, nc26585, nc26586, dw[21]}),
		.dipa (),
		.dipb (),
		.cea (net_592),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_332 (
		.doa ({nc26587, nc26588, nc26589, nc26590, nc26591, nc26592, nc26593, nc26594, nc26595, nc26596, nc26597, nc26598, nc26599, nc26600, nc26601, nc26602, nc26603, nc26604, nc26605, nc26606, nc26607, nc26608, nc26609, nc26610, nc26611, nc26612, nc26613, nc26614, nc26615, nc26616, nc26617, nc26618, nc26619, nc26620, nc26621, nc26622, nc26623, nc26624, nc26625, nc26626, nc26627, nc26628, nc26629, nc26630, nc26631, nc26632, nc26633, nc26634, nc26635, nc26636, nc26637, nc26638, nc26639, nc26640, nc26641, nc26642, nc26643, nc26644, nc26645, nc26646, nc26647, nc26648, nc26649, net_598}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26650, nc26651, nc26652, nc26653, nc26654, nc26655, nc26656, nc26657, nc26658, nc26659, nc26660, nc26661, nc26662, nc26663, nc26664, nc26665, nc26666, nc26667, nc26668, nc26669, nc26670, nc26671, nc26672, nc26673, nc26674, nc26675, nc26676, nc26677, nc26678, nc26679, nc26680, nc26681, nc26682, nc26683, nc26684, nc26685, nc26686, nc26687, nc26688, nc26689, nc26690, nc26691, nc26692, nc26693, nc26694, nc26695, nc26696, nc26697, nc26698, nc26699, nc26700, nc26701, nc26702, nc26703, nc26704, nc26705, nc26706, nc26707, nc26708, nc26709, nc26710, nc26711, nc26712, dw[29]}),
		.dipa (),
		.dipb (),
		.cea (net_596),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u304 (
		.sel (addra_pipe_0_net),
		.i0 (net_594),
		.i1 (net_598),
		.o (net_600)
	);
fifo2ram_emb_v1_AND u305 (
		.i0 (net_602),
		.i1 (net_601),
		.o (net_592)
	);
fifo2ram_emb_v1_AND u306 (
		.i0 (net_602),
		.i1 (ar[0]),
		.o (net_596)
	);
fifo2ram_emb_v1_NOT u307 (
		.i (ar[0]),
		.o (net_601)
	);
fifo2ram_emb_v1_MUX u308 (
		.sel (addra_pipe_1_net),
		.i0 (net_589),
		.i1 (net_600),
		.o (net_603)
	);
fifo2ram_emb_v1_AND u309 (
		.i0 (net_605),
		.i1 (net_604),
		.o (net_591)
	);
fifo2ram_emb_v1_AND u310 (
		.i0 (net_605),
		.i1 (ar[1]),
		.o (net_602)
	);
fifo2ram_emb_v1_NOT u311 (
		.i (ar[1]),
		.o (net_604)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_336 (
		.doa ({nc26713, nc26714, nc26715, nc26716, nc26717, nc26718, nc26719, nc26720, nc26721, nc26722, nc26723, nc26724, nc26725, nc26726, nc26727, nc26728, nc26729, nc26730, nc26731, nc26732, nc26733, nc26734, nc26735, nc26736, nc26737, nc26738, nc26739, nc26740, nc26741, nc26742, nc26743, nc26744, nc26745, nc26746, nc26747, nc26748, nc26749, nc26750, nc26751, nc26752, nc26753, nc26754, nc26755, nc26756, nc26757, nc26758, nc26759, nc26760, nc26761, nc26762, nc26763, nc26764, nc26765, nc26766, nc26767, nc26768, nc26769, nc26770, nc26771, nc26772, nc26773, nc26774, nc26775, net_608}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26776, nc26777, nc26778, nc26779, nc26780, nc26781, nc26782, nc26783, nc26784, nc26785, nc26786, nc26787, nc26788, nc26789, nc26790, nc26791, nc26792, nc26793, nc26794, nc26795, nc26796, nc26797, nc26798, nc26799, nc26800, nc26801, nc26802, nc26803, nc26804, nc26805, nc26806, nc26807, nc26808, nc26809, nc26810, nc26811, nc26812, nc26813, nc26814, nc26815, nc26816, nc26817, nc26818, nc26819, nc26820, nc26821, nc26822, nc26823, nc26824, nc26825, nc26826, nc26827, nc26828, nc26829, nc26830, nc26831, nc26832, nc26833, nc26834, nc26835, nc26836, nc26837, nc26838, dw[37]}),
		.dipa (),
		.dipb (),
		.cea (net_606),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_340 (
		.doa ({nc26839, nc26840, nc26841, nc26842, nc26843, nc26844, nc26845, nc26846, nc26847, nc26848, nc26849, nc26850, nc26851, nc26852, nc26853, nc26854, nc26855, nc26856, nc26857, nc26858, nc26859, nc26860, nc26861, nc26862, nc26863, nc26864, nc26865, nc26866, nc26867, nc26868, nc26869, nc26870, nc26871, nc26872, nc26873, nc26874, nc26875, nc26876, nc26877, nc26878, nc26879, nc26880, nc26881, nc26882, nc26883, nc26884, nc26885, nc26886, nc26887, nc26888, nc26889, nc26890, nc26891, nc26892, nc26893, nc26894, nc26895, nc26896, nc26897, nc26898, nc26899, nc26900, nc26901, net_612}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc26902, nc26903, nc26904, nc26905, nc26906, nc26907, nc26908, nc26909, nc26910, nc26911, nc26912, nc26913, nc26914, nc26915, nc26916, nc26917, nc26918, nc26919, nc26920, nc26921, nc26922, nc26923, nc26924, nc26925, nc26926, nc26927, nc26928, nc26929, nc26930, nc26931, nc26932, nc26933, nc26934, nc26935, nc26936, nc26937, nc26938, nc26939, nc26940, nc26941, nc26942, nc26943, nc26944, nc26945, nc26946, nc26947, nc26948, nc26949, nc26950, nc26951, nc26952, nc26953, nc26954, nc26955, nc26956, nc26957, nc26958, nc26959, nc26960, nc26961, nc26962, nc26963, nc26964, dw[45]}),
		.dipa (),
		.dipb (),
		.cea (net_610),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u312 (
		.sel (addra_pipe_0_net),
		.i0 (net_608),
		.i1 (net_612),
		.o (net_614)
	);
fifo2ram_emb_v1_AND u313 (
		.i0 (net_616),
		.i1 (net_615),
		.o (net_606)
	);
fifo2ram_emb_v1_AND u314 (
		.i0 (net_616),
		.i1 (ar[0]),
		.o (net_610)
	);
fifo2ram_emb_v1_NOT u315 (
		.i (ar[0]),
		.o (net_615)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_344 (
		.doa ({nc26965, nc26966, nc26967, nc26968, nc26969, nc26970, nc26971, nc26972, nc26973, nc26974, nc26975, nc26976, nc26977, nc26978, nc26979, nc26980, nc26981, nc26982, nc26983, nc26984, nc26985, nc26986, nc26987, nc26988, nc26989, nc26990, nc26991, nc26992, nc26993, nc26994, nc26995, nc26996, nc26997, nc26998, nc26999, nc27000, nc27001, nc27002, nc27003, nc27004, nc27005, nc27006, nc27007, nc27008, nc27009, nc27010, nc27011, nc27012, nc27013, nc27014, nc27015, nc27016, nc27017, nc27018, nc27019, nc27020, nc27021, nc27022, nc27023, nc27024, nc27025, nc27026, nc27027, net_619}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27028, nc27029, nc27030, nc27031, nc27032, nc27033, nc27034, nc27035, nc27036, nc27037, nc27038, nc27039, nc27040, nc27041, nc27042, nc27043, nc27044, nc27045, nc27046, nc27047, nc27048, nc27049, nc27050, nc27051, nc27052, nc27053, nc27054, nc27055, nc27056, nc27057, nc27058, nc27059, nc27060, nc27061, nc27062, nc27063, nc27064, nc27065, nc27066, nc27067, nc27068, nc27069, nc27070, nc27071, nc27072, nc27073, nc27074, nc27075, nc27076, nc27077, nc27078, nc27079, nc27080, nc27081, nc27082, nc27083, nc27084, nc27085, nc27086, nc27087, nc27088, nc27089, nc27090, dw[53]}),
		.dipa (),
		.dipb (),
		.cea (net_617),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_348 (
		.doa ({nc27091, nc27092, nc27093, nc27094, nc27095, nc27096, nc27097, nc27098, nc27099, nc27100, nc27101, nc27102, nc27103, nc27104, nc27105, nc27106, nc27107, nc27108, nc27109, nc27110, nc27111, nc27112, nc27113, nc27114, nc27115, nc27116, nc27117, nc27118, nc27119, nc27120, nc27121, nc27122, nc27123, nc27124, nc27125, nc27126, nc27127, nc27128, nc27129, nc27130, nc27131, nc27132, nc27133, nc27134, nc27135, nc27136, nc27137, nc27138, nc27139, nc27140, nc27141, nc27142, nc27143, nc27144, nc27145, nc27146, nc27147, nc27148, nc27149, nc27150, nc27151, nc27152, nc27153, net_623}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27154, nc27155, nc27156, nc27157, nc27158, nc27159, nc27160, nc27161, nc27162, nc27163, nc27164, nc27165, nc27166, nc27167, nc27168, nc27169, nc27170, nc27171, nc27172, nc27173, nc27174, nc27175, nc27176, nc27177, nc27178, nc27179, nc27180, nc27181, nc27182, nc27183, nc27184, nc27185, nc27186, nc27187, nc27188, nc27189, nc27190, nc27191, nc27192, nc27193, nc27194, nc27195, nc27196, nc27197, nc27198, nc27199, nc27200, nc27201, nc27202, nc27203, nc27204, nc27205, nc27206, nc27207, nc27208, nc27209, nc27210, nc27211, nc27212, nc27213, nc27214, nc27215, nc27216, dw[61]}),
		.dipa (),
		.dipb (),
		.cea (net_621),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u316 (
		.sel (addra_pipe_0_net),
		.i0 (net_619),
		.i1 (net_623),
		.o (net_625)
	);
fifo2ram_emb_v1_AND u317 (
		.i0 (net_627),
		.i1 (net_626),
		.o (net_617)
	);
fifo2ram_emb_v1_AND u318 (
		.i0 (net_627),
		.i1 (ar[0]),
		.o (net_621)
	);
fifo2ram_emb_v1_NOT u319 (
		.i (ar[0]),
		.o (net_626)
	);
fifo2ram_emb_v1_MUX u320 (
		.sel (addra_pipe_1_net),
		.i0 (net_614),
		.i1 (net_625),
		.o (net_628)
	);
fifo2ram_emb_v1_AND u321 (
		.i0 (net_630),
		.i1 (net_629),
		.o (net_616)
	);
fifo2ram_emb_v1_AND u322 (
		.i0 (net_630),
		.i1 (ar[1]),
		.o (net_627)
	);
fifo2ram_emb_v1_NOT u323 (
		.i (ar[1]),
		.o (net_629)
	);
fifo2ram_emb_v1_MUX u324 (
		.sel (addra_pipe_2_net),
		.i0 (net_603),
		.i1 (net_628),
		.o (net_631)
	);
fifo2ram_emb_v1_AND u325 (
		.i0 (net_633),
		.i1 (net_632),
		.o (net_605)
	);
fifo2ram_emb_v1_AND u326 (
		.i0 (net_633),
		.i1 (ar[2]),
		.o (net_630)
	);
fifo2ram_emb_v1_NOT u327 (
		.i (ar[2]),
		.o (net_632)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_352 (
		.doa ({nc27217, nc27218, nc27219, nc27220, nc27221, nc27222, nc27223, nc27224, nc27225, nc27226, nc27227, nc27228, nc27229, nc27230, nc27231, nc27232, nc27233, nc27234, nc27235, nc27236, nc27237, nc27238, nc27239, nc27240, nc27241, nc27242, nc27243, nc27244, nc27245, nc27246, nc27247, nc27248, nc27249, nc27250, nc27251, nc27252, nc27253, nc27254, nc27255, nc27256, nc27257, nc27258, nc27259, nc27260, nc27261, nc27262, nc27263, nc27264, nc27265, nc27266, nc27267, nc27268, nc27269, nc27270, nc27271, nc27272, nc27273, nc27274, nc27275, nc27276, nc27277, nc27278, nc27279, net_636}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27280, nc27281, nc27282, nc27283, nc27284, nc27285, nc27286, nc27287, nc27288, nc27289, nc27290, nc27291, nc27292, nc27293, nc27294, nc27295, nc27296, nc27297, nc27298, nc27299, nc27300, nc27301, nc27302, nc27303, nc27304, nc27305, nc27306, nc27307, nc27308, nc27309, nc27310, nc27311, nc27312, nc27313, nc27314, nc27315, nc27316, nc27317, nc27318, nc27319, nc27320, nc27321, nc27322, nc27323, nc27324, nc27325, nc27326, nc27327, nc27328, nc27329, nc27330, nc27331, nc27332, nc27333, nc27334, nc27335, nc27336, nc27337, nc27338, nc27339, nc27340, nc27341, nc27342, dw[69]}),
		.dipa (),
		.dipb (),
		.cea (net_634),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_356 (
		.doa ({nc27343, nc27344, nc27345, nc27346, nc27347, nc27348, nc27349, nc27350, nc27351, nc27352, nc27353, nc27354, nc27355, nc27356, nc27357, nc27358, nc27359, nc27360, nc27361, nc27362, nc27363, nc27364, nc27365, nc27366, nc27367, nc27368, nc27369, nc27370, nc27371, nc27372, nc27373, nc27374, nc27375, nc27376, nc27377, nc27378, nc27379, nc27380, nc27381, nc27382, nc27383, nc27384, nc27385, nc27386, nc27387, nc27388, nc27389, nc27390, nc27391, nc27392, nc27393, nc27394, nc27395, nc27396, nc27397, nc27398, nc27399, nc27400, nc27401, nc27402, nc27403, nc27404, nc27405, net_640}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27406, nc27407, nc27408, nc27409, nc27410, nc27411, nc27412, nc27413, nc27414, nc27415, nc27416, nc27417, nc27418, nc27419, nc27420, nc27421, nc27422, nc27423, nc27424, nc27425, nc27426, nc27427, nc27428, nc27429, nc27430, nc27431, nc27432, nc27433, nc27434, nc27435, nc27436, nc27437, nc27438, nc27439, nc27440, nc27441, nc27442, nc27443, nc27444, nc27445, nc27446, nc27447, nc27448, nc27449, nc27450, nc27451, nc27452, nc27453, nc27454, nc27455, nc27456, nc27457, nc27458, nc27459, nc27460, nc27461, nc27462, nc27463, nc27464, nc27465, nc27466, nc27467, nc27468, dw[77]}),
		.dipa (),
		.dipb (),
		.cea (net_638),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u328 (
		.sel (addra_pipe_0_net),
		.i0 (net_636),
		.i1 (net_640),
		.o (net_642)
	);
fifo2ram_emb_v1_AND u329 (
		.i0 (net_644),
		.i1 (net_643),
		.o (net_634)
	);
fifo2ram_emb_v1_AND u330 (
		.i0 (net_644),
		.i1 (ar[0]),
		.o (net_638)
	);
fifo2ram_emb_v1_NOT u331 (
		.i (ar[0]),
		.o (net_643)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_360 (
		.doa ({nc27469, nc27470, nc27471, nc27472, nc27473, nc27474, nc27475, nc27476, nc27477, nc27478, nc27479, nc27480, nc27481, nc27482, nc27483, nc27484, nc27485, nc27486, nc27487, nc27488, nc27489, nc27490, nc27491, nc27492, nc27493, nc27494, nc27495, nc27496, nc27497, nc27498, nc27499, nc27500, nc27501, nc27502, nc27503, nc27504, nc27505, nc27506, nc27507, nc27508, nc27509, nc27510, nc27511, nc27512, nc27513, nc27514, nc27515, nc27516, nc27517, nc27518, nc27519, nc27520, nc27521, nc27522, nc27523, nc27524, nc27525, nc27526, nc27527, nc27528, nc27529, nc27530, nc27531, net_647}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27532, nc27533, nc27534, nc27535, nc27536, nc27537, nc27538, nc27539, nc27540, nc27541, nc27542, nc27543, nc27544, nc27545, nc27546, nc27547, nc27548, nc27549, nc27550, nc27551, nc27552, nc27553, nc27554, nc27555, nc27556, nc27557, nc27558, nc27559, nc27560, nc27561, nc27562, nc27563, nc27564, nc27565, nc27566, nc27567, nc27568, nc27569, nc27570, nc27571, nc27572, nc27573, nc27574, nc27575, nc27576, nc27577, nc27578, nc27579, nc27580, nc27581, nc27582, nc27583, nc27584, nc27585, nc27586, nc27587, nc27588, nc27589, nc27590, nc27591, nc27592, nc27593, nc27594, dw[85]}),
		.dipa (),
		.dipb (),
		.cea (net_645),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_364 (
		.doa ({nc27595, nc27596, nc27597, nc27598, nc27599, nc27600, nc27601, nc27602, nc27603, nc27604, nc27605, nc27606, nc27607, nc27608, nc27609, nc27610, nc27611, nc27612, nc27613, nc27614, nc27615, nc27616, nc27617, nc27618, nc27619, nc27620, nc27621, nc27622, nc27623, nc27624, nc27625, nc27626, nc27627, nc27628, nc27629, nc27630, nc27631, nc27632, nc27633, nc27634, nc27635, nc27636, nc27637, nc27638, nc27639, nc27640, nc27641, nc27642, nc27643, nc27644, nc27645, nc27646, nc27647, nc27648, nc27649, nc27650, nc27651, nc27652, nc27653, nc27654, nc27655, nc27656, nc27657, net_651}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27658, nc27659, nc27660, nc27661, nc27662, nc27663, nc27664, nc27665, nc27666, nc27667, nc27668, nc27669, nc27670, nc27671, nc27672, nc27673, nc27674, nc27675, nc27676, nc27677, nc27678, nc27679, nc27680, nc27681, nc27682, nc27683, nc27684, nc27685, nc27686, nc27687, nc27688, nc27689, nc27690, nc27691, nc27692, nc27693, nc27694, nc27695, nc27696, nc27697, nc27698, nc27699, nc27700, nc27701, nc27702, nc27703, nc27704, nc27705, nc27706, nc27707, nc27708, nc27709, nc27710, nc27711, nc27712, nc27713, nc27714, nc27715, nc27716, nc27717, nc27718, nc27719, nc27720, dw[93]}),
		.dipa (),
		.dipb (),
		.cea (net_649),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u332 (
		.sel (addra_pipe_0_net),
		.i0 (net_647),
		.i1 (net_651),
		.o (net_653)
	);
fifo2ram_emb_v1_AND u333 (
		.i0 (net_655),
		.i1 (net_654),
		.o (net_645)
	);
fifo2ram_emb_v1_AND u334 (
		.i0 (net_655),
		.i1 (ar[0]),
		.o (net_649)
	);
fifo2ram_emb_v1_NOT u335 (
		.i (ar[0]),
		.o (net_654)
	);
fifo2ram_emb_v1_MUX u336 (
		.sel (addra_pipe_1_net),
		.i0 (net_642),
		.i1 (net_653),
		.o (net_656)
	);
fifo2ram_emb_v1_AND u337 (
		.i0 (net_658),
		.i1 (net_657),
		.o (net_644)
	);
fifo2ram_emb_v1_AND u338 (
		.i0 (net_658),
		.i1 (ar[1]),
		.o (net_655)
	);
fifo2ram_emb_v1_NOT u339 (
		.i (ar[1]),
		.o (net_657)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_368 (
		.doa ({nc27721, nc27722, nc27723, nc27724, nc27725, nc27726, nc27727, nc27728, nc27729, nc27730, nc27731, nc27732, nc27733, nc27734, nc27735, nc27736, nc27737, nc27738, nc27739, nc27740, nc27741, nc27742, nc27743, nc27744, nc27745, nc27746, nc27747, nc27748, nc27749, nc27750, nc27751, nc27752, nc27753, nc27754, nc27755, nc27756, nc27757, nc27758, nc27759, nc27760, nc27761, nc27762, nc27763, nc27764, nc27765, nc27766, nc27767, nc27768, nc27769, nc27770, nc27771, nc27772, nc27773, nc27774, nc27775, nc27776, nc27777, nc27778, nc27779, nc27780, nc27781, nc27782, nc27783, net_661}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27784, nc27785, nc27786, nc27787, nc27788, nc27789, nc27790, nc27791, nc27792, nc27793, nc27794, nc27795, nc27796, nc27797, nc27798, nc27799, nc27800, nc27801, nc27802, nc27803, nc27804, nc27805, nc27806, nc27807, nc27808, nc27809, nc27810, nc27811, nc27812, nc27813, nc27814, nc27815, nc27816, nc27817, nc27818, nc27819, nc27820, nc27821, nc27822, nc27823, nc27824, nc27825, nc27826, nc27827, nc27828, nc27829, nc27830, nc27831, nc27832, nc27833, nc27834, nc27835, nc27836, nc27837, nc27838, nc27839, nc27840, nc27841, nc27842, nc27843, nc27844, nc27845, nc27846, dw[101]}),
		.dipa (),
		.dipb (),
		.cea (net_659),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_372 (
		.doa ({nc27847, nc27848, nc27849, nc27850, nc27851, nc27852, nc27853, nc27854, nc27855, nc27856, nc27857, nc27858, nc27859, nc27860, nc27861, nc27862, nc27863, nc27864, nc27865, nc27866, nc27867, nc27868, nc27869, nc27870, nc27871, nc27872, nc27873, nc27874, nc27875, nc27876, nc27877, nc27878, nc27879, nc27880, nc27881, nc27882, nc27883, nc27884, nc27885, nc27886, nc27887, nc27888, nc27889, nc27890, nc27891, nc27892, nc27893, nc27894, nc27895, nc27896, nc27897, nc27898, nc27899, nc27900, nc27901, nc27902, nc27903, nc27904, nc27905, nc27906, nc27907, nc27908, nc27909, net_665}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc27910, nc27911, nc27912, nc27913, nc27914, nc27915, nc27916, nc27917, nc27918, nc27919, nc27920, nc27921, nc27922, nc27923, nc27924, nc27925, nc27926, nc27927, nc27928, nc27929, nc27930, nc27931, nc27932, nc27933, nc27934, nc27935, nc27936, nc27937, nc27938, nc27939, nc27940, nc27941, nc27942, nc27943, nc27944, nc27945, nc27946, nc27947, nc27948, nc27949, nc27950, nc27951, nc27952, nc27953, nc27954, nc27955, nc27956, nc27957, nc27958, nc27959, nc27960, nc27961, nc27962, nc27963, nc27964, nc27965, nc27966, nc27967, nc27968, nc27969, nc27970, nc27971, nc27972, dw[109]}),
		.dipa (),
		.dipb (),
		.cea (net_663),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u340 (
		.sel (addra_pipe_0_net),
		.i0 (net_661),
		.i1 (net_665),
		.o (net_667)
	);
fifo2ram_emb_v1_AND u341 (
		.i0 (net_669),
		.i1 (net_668),
		.o (net_659)
	);
fifo2ram_emb_v1_AND u342 (
		.i0 (net_669),
		.i1 (ar[0]),
		.o (net_663)
	);
fifo2ram_emb_v1_NOT u343 (
		.i (ar[0]),
		.o (net_668)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_376 (
		.doa ({nc27973, nc27974, nc27975, nc27976, nc27977, nc27978, nc27979, nc27980, nc27981, nc27982, nc27983, nc27984, nc27985, nc27986, nc27987, nc27988, nc27989, nc27990, nc27991, nc27992, nc27993, nc27994, nc27995, nc27996, nc27997, nc27998, nc27999, nc28000, nc28001, nc28002, nc28003, nc28004, nc28005, nc28006, nc28007, nc28008, nc28009, nc28010, nc28011, nc28012, nc28013, nc28014, nc28015, nc28016, nc28017, nc28018, nc28019, nc28020, nc28021, nc28022, nc28023, nc28024, nc28025, nc28026, nc28027, nc28028, nc28029, nc28030, nc28031, nc28032, nc28033, nc28034, nc28035, net_672}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28036, nc28037, nc28038, nc28039, nc28040, nc28041, nc28042, nc28043, nc28044, nc28045, nc28046, nc28047, nc28048, nc28049, nc28050, nc28051, nc28052, nc28053, nc28054, nc28055, nc28056, nc28057, nc28058, nc28059, nc28060, nc28061, nc28062, nc28063, nc28064, nc28065, nc28066, nc28067, nc28068, nc28069, nc28070, nc28071, nc28072, nc28073, nc28074, nc28075, nc28076, nc28077, nc28078, nc28079, nc28080, nc28081, nc28082, nc28083, nc28084, nc28085, nc28086, nc28087, nc28088, nc28089, nc28090, nc28091, nc28092, nc28093, nc28094, nc28095, nc28096, nc28097, nc28098, dw[117]}),
		.dipa (),
		.dipb (),
		.cea (net_670),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_380 (
		.doa ({nc28099, nc28100, nc28101, nc28102, nc28103, nc28104, nc28105, nc28106, nc28107, nc28108, nc28109, nc28110, nc28111, nc28112, nc28113, nc28114, nc28115, nc28116, nc28117, nc28118, nc28119, nc28120, nc28121, nc28122, nc28123, nc28124, nc28125, nc28126, nc28127, nc28128, nc28129, nc28130, nc28131, nc28132, nc28133, nc28134, nc28135, nc28136, nc28137, nc28138, nc28139, nc28140, nc28141, nc28142, nc28143, nc28144, nc28145, nc28146, nc28147, nc28148, nc28149, nc28150, nc28151, nc28152, nc28153, nc28154, nc28155, nc28156, nc28157, nc28158, nc28159, nc28160, nc28161, net_676}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28162, nc28163, nc28164, nc28165, nc28166, nc28167, nc28168, nc28169, nc28170, nc28171, nc28172, nc28173, nc28174, nc28175, nc28176, nc28177, nc28178, nc28179, nc28180, nc28181, nc28182, nc28183, nc28184, nc28185, nc28186, nc28187, nc28188, nc28189, nc28190, nc28191, nc28192, nc28193, nc28194, nc28195, nc28196, nc28197, nc28198, nc28199, nc28200, nc28201, nc28202, nc28203, nc28204, nc28205, nc28206, nc28207, nc28208, nc28209, nc28210, nc28211, nc28212, nc28213, nc28214, nc28215, nc28216, nc28217, nc28218, nc28219, nc28220, nc28221, nc28222, nc28223, nc28224, dw[125]}),
		.dipa (),
		.dipb (),
		.cea (net_674),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u344 (
		.sel (addra_pipe_0_net),
		.i0 (net_672),
		.i1 (net_676),
		.o (net_678)
	);
fifo2ram_emb_v1_AND u345 (
		.i0 (net_680),
		.i1 (net_679),
		.o (net_670)
	);
fifo2ram_emb_v1_AND u346 (
		.i0 (net_680),
		.i1 (ar[0]),
		.o (net_674)
	);
fifo2ram_emb_v1_NOT u347 (
		.i (ar[0]),
		.o (net_679)
	);
fifo2ram_emb_v1_MUX u348 (
		.sel (addra_pipe_1_net),
		.i0 (net_667),
		.i1 (net_678),
		.o (net_681)
	);
fifo2ram_emb_v1_AND u349 (
		.i0 (net_683),
		.i1 (net_682),
		.o (net_669)
	);
fifo2ram_emb_v1_AND u350 (
		.i0 (net_683),
		.i1 (ar[1]),
		.o (net_680)
	);
fifo2ram_emb_v1_NOT u351 (
		.i (ar[1]),
		.o (net_682)
	);
fifo2ram_emb_v1_MUX u352 (
		.sel (addra_pipe_2_net),
		.i0 (net_656),
		.i1 (net_681),
		.o (net_684)
	);
fifo2ram_emb_v1_AND u353 (
		.i0 (net_686),
		.i1 (net_685),
		.o (net_658)
	);
fifo2ram_emb_v1_AND u354 (
		.i0 (net_686),
		.i1 (ar[2]),
		.o (net_683)
	);
fifo2ram_emb_v1_NOT u355 (
		.i (ar[2]),
		.o (net_685)
	);
fifo2ram_emb_v1_MUX u356 (
		.sel (addra_pipe_3_net),
		.i0 (net_631),
		.i1 (net_684),
		.o (qr[5])
	);
fifo2ram_emb_v1_AND u357 (
		.i0 (cer),
		.i1 (net_688),
		.o (net_633)
	);
fifo2ram_emb_v1_AND u358 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_686)
	);
fifo2ram_emb_v1_NOT u359 (
		.i (ar[3]),
		.o (net_688)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_384 (
		.doa ({nc28225, nc28226, nc28227, nc28228, nc28229, nc28230, nc28231, nc28232, nc28233, nc28234, nc28235, nc28236, nc28237, nc28238, nc28239, nc28240, nc28241, nc28242, nc28243, nc28244, nc28245, nc28246, nc28247, nc28248, nc28249, nc28250, nc28251, nc28252, nc28253, nc28254, nc28255, nc28256, nc28257, nc28258, nc28259, nc28260, nc28261, nc28262, nc28263, nc28264, nc28265, nc28266, nc28267, nc28268, nc28269, nc28270, nc28271, nc28272, nc28273, nc28274, nc28275, nc28276, nc28277, nc28278, nc28279, nc28280, nc28281, nc28282, nc28283, nc28284, nc28285, nc28286, nc28287, net_692}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28288, nc28289, nc28290, nc28291, nc28292, nc28293, nc28294, nc28295, nc28296, nc28297, nc28298, nc28299, nc28300, nc28301, nc28302, nc28303, nc28304, nc28305, nc28306, nc28307, nc28308, nc28309, nc28310, nc28311, nc28312, nc28313, nc28314, nc28315, nc28316, nc28317, nc28318, nc28319, nc28320, nc28321, nc28322, nc28323, nc28324, nc28325, nc28326, nc28327, nc28328, nc28329, nc28330, nc28331, nc28332, nc28333, nc28334, nc28335, nc28336, nc28337, nc28338, nc28339, nc28340, nc28341, nc28342, nc28343, nc28344, nc28345, nc28346, nc28347, nc28348, nc28349, nc28350, dw[6]}),
		.dipa (),
		.dipb (),
		.cea (net_690),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_388 (
		.doa ({nc28351, nc28352, nc28353, nc28354, nc28355, nc28356, nc28357, nc28358, nc28359, nc28360, nc28361, nc28362, nc28363, nc28364, nc28365, nc28366, nc28367, nc28368, nc28369, nc28370, nc28371, nc28372, nc28373, nc28374, nc28375, nc28376, nc28377, nc28378, nc28379, nc28380, nc28381, nc28382, nc28383, nc28384, nc28385, nc28386, nc28387, nc28388, nc28389, nc28390, nc28391, nc28392, nc28393, nc28394, nc28395, nc28396, nc28397, nc28398, nc28399, nc28400, nc28401, nc28402, nc28403, nc28404, nc28405, nc28406, nc28407, nc28408, nc28409, nc28410, nc28411, nc28412, nc28413, net_696}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28414, nc28415, nc28416, nc28417, nc28418, nc28419, nc28420, nc28421, nc28422, nc28423, nc28424, nc28425, nc28426, nc28427, nc28428, nc28429, nc28430, nc28431, nc28432, nc28433, nc28434, nc28435, nc28436, nc28437, nc28438, nc28439, nc28440, nc28441, nc28442, nc28443, nc28444, nc28445, nc28446, nc28447, nc28448, nc28449, nc28450, nc28451, nc28452, nc28453, nc28454, nc28455, nc28456, nc28457, nc28458, nc28459, nc28460, nc28461, nc28462, nc28463, nc28464, nc28465, nc28466, nc28467, nc28468, nc28469, nc28470, nc28471, nc28472, nc28473, nc28474, nc28475, nc28476, dw[14]}),
		.dipa (),
		.dipb (),
		.cea (net_694),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u360 (
		.sel (addra_pipe_0_net),
		.i0 (net_692),
		.i1 (net_696),
		.o (net_698)
	);
fifo2ram_emb_v1_AND u361 (
		.i0 (net_700),
		.i1 (net_699),
		.o (net_690)
	);
fifo2ram_emb_v1_AND u362 (
		.i0 (net_700),
		.i1 (ar[0]),
		.o (net_694)
	);
fifo2ram_emb_v1_NOT u363 (
		.i (ar[0]),
		.o (net_699)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_392 (
		.doa ({nc28477, nc28478, nc28479, nc28480, nc28481, nc28482, nc28483, nc28484, nc28485, nc28486, nc28487, nc28488, nc28489, nc28490, nc28491, nc28492, nc28493, nc28494, nc28495, nc28496, nc28497, nc28498, nc28499, nc28500, nc28501, nc28502, nc28503, nc28504, nc28505, nc28506, nc28507, nc28508, nc28509, nc28510, nc28511, nc28512, nc28513, nc28514, nc28515, nc28516, nc28517, nc28518, nc28519, nc28520, nc28521, nc28522, nc28523, nc28524, nc28525, nc28526, nc28527, nc28528, nc28529, nc28530, nc28531, nc28532, nc28533, nc28534, nc28535, nc28536, nc28537, nc28538, nc28539, net_703}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28540, nc28541, nc28542, nc28543, nc28544, nc28545, nc28546, nc28547, nc28548, nc28549, nc28550, nc28551, nc28552, nc28553, nc28554, nc28555, nc28556, nc28557, nc28558, nc28559, nc28560, nc28561, nc28562, nc28563, nc28564, nc28565, nc28566, nc28567, nc28568, nc28569, nc28570, nc28571, nc28572, nc28573, nc28574, nc28575, nc28576, nc28577, nc28578, nc28579, nc28580, nc28581, nc28582, nc28583, nc28584, nc28585, nc28586, nc28587, nc28588, nc28589, nc28590, nc28591, nc28592, nc28593, nc28594, nc28595, nc28596, nc28597, nc28598, nc28599, nc28600, nc28601, nc28602, dw[22]}),
		.dipa (),
		.dipb (),
		.cea (net_701),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_396 (
		.doa ({nc28603, nc28604, nc28605, nc28606, nc28607, nc28608, nc28609, nc28610, nc28611, nc28612, nc28613, nc28614, nc28615, nc28616, nc28617, nc28618, nc28619, nc28620, nc28621, nc28622, nc28623, nc28624, nc28625, nc28626, nc28627, nc28628, nc28629, nc28630, nc28631, nc28632, nc28633, nc28634, nc28635, nc28636, nc28637, nc28638, nc28639, nc28640, nc28641, nc28642, nc28643, nc28644, nc28645, nc28646, nc28647, nc28648, nc28649, nc28650, nc28651, nc28652, nc28653, nc28654, nc28655, nc28656, nc28657, nc28658, nc28659, nc28660, nc28661, nc28662, nc28663, nc28664, nc28665, net_707}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28666, nc28667, nc28668, nc28669, nc28670, nc28671, nc28672, nc28673, nc28674, nc28675, nc28676, nc28677, nc28678, nc28679, nc28680, nc28681, nc28682, nc28683, nc28684, nc28685, nc28686, nc28687, nc28688, nc28689, nc28690, nc28691, nc28692, nc28693, nc28694, nc28695, nc28696, nc28697, nc28698, nc28699, nc28700, nc28701, nc28702, nc28703, nc28704, nc28705, nc28706, nc28707, nc28708, nc28709, nc28710, nc28711, nc28712, nc28713, nc28714, nc28715, nc28716, nc28717, nc28718, nc28719, nc28720, nc28721, nc28722, nc28723, nc28724, nc28725, nc28726, nc28727, nc28728, dw[30]}),
		.dipa (),
		.dipb (),
		.cea (net_705),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u364 (
		.sel (addra_pipe_0_net),
		.i0 (net_703),
		.i1 (net_707),
		.o (net_709)
	);
fifo2ram_emb_v1_AND u365 (
		.i0 (net_711),
		.i1 (net_710),
		.o (net_701)
	);
fifo2ram_emb_v1_AND u366 (
		.i0 (net_711),
		.i1 (ar[0]),
		.o (net_705)
	);
fifo2ram_emb_v1_NOT u367 (
		.i (ar[0]),
		.o (net_710)
	);
fifo2ram_emb_v1_MUX u368 (
		.sel (addra_pipe_1_net),
		.i0 (net_698),
		.i1 (net_709),
		.o (net_712)
	);
fifo2ram_emb_v1_AND u369 (
		.i0 (net_714),
		.i1 (net_713),
		.o (net_700)
	);
fifo2ram_emb_v1_AND u370 (
		.i0 (net_714),
		.i1 (ar[1]),
		.o (net_711)
	);
fifo2ram_emb_v1_NOT u371 (
		.i (ar[1]),
		.o (net_713)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_400 (
		.doa ({nc28729, nc28730, nc28731, nc28732, nc28733, nc28734, nc28735, nc28736, nc28737, nc28738, nc28739, nc28740, nc28741, nc28742, nc28743, nc28744, nc28745, nc28746, nc28747, nc28748, nc28749, nc28750, nc28751, nc28752, nc28753, nc28754, nc28755, nc28756, nc28757, nc28758, nc28759, nc28760, nc28761, nc28762, nc28763, nc28764, nc28765, nc28766, nc28767, nc28768, nc28769, nc28770, nc28771, nc28772, nc28773, nc28774, nc28775, nc28776, nc28777, nc28778, nc28779, nc28780, nc28781, nc28782, nc28783, nc28784, nc28785, nc28786, nc28787, nc28788, nc28789, nc28790, nc28791, net_717}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28792, nc28793, nc28794, nc28795, nc28796, nc28797, nc28798, nc28799, nc28800, nc28801, nc28802, nc28803, nc28804, nc28805, nc28806, nc28807, nc28808, nc28809, nc28810, nc28811, nc28812, nc28813, nc28814, nc28815, nc28816, nc28817, nc28818, nc28819, nc28820, nc28821, nc28822, nc28823, nc28824, nc28825, nc28826, nc28827, nc28828, nc28829, nc28830, nc28831, nc28832, nc28833, nc28834, nc28835, nc28836, nc28837, nc28838, nc28839, nc28840, nc28841, nc28842, nc28843, nc28844, nc28845, nc28846, nc28847, nc28848, nc28849, nc28850, nc28851, nc28852, nc28853, nc28854, dw[38]}),
		.dipa (),
		.dipb (),
		.cea (net_715),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_404 (
		.doa ({nc28855, nc28856, nc28857, nc28858, nc28859, nc28860, nc28861, nc28862, nc28863, nc28864, nc28865, nc28866, nc28867, nc28868, nc28869, nc28870, nc28871, nc28872, nc28873, nc28874, nc28875, nc28876, nc28877, nc28878, nc28879, nc28880, nc28881, nc28882, nc28883, nc28884, nc28885, nc28886, nc28887, nc28888, nc28889, nc28890, nc28891, nc28892, nc28893, nc28894, nc28895, nc28896, nc28897, nc28898, nc28899, nc28900, nc28901, nc28902, nc28903, nc28904, nc28905, nc28906, nc28907, nc28908, nc28909, nc28910, nc28911, nc28912, nc28913, nc28914, nc28915, nc28916, nc28917, net_721}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc28918, nc28919, nc28920, nc28921, nc28922, nc28923, nc28924, nc28925, nc28926, nc28927, nc28928, nc28929, nc28930, nc28931, nc28932, nc28933, nc28934, nc28935, nc28936, nc28937, nc28938, nc28939, nc28940, nc28941, nc28942, nc28943, nc28944, nc28945, nc28946, nc28947, nc28948, nc28949, nc28950, nc28951, nc28952, nc28953, nc28954, nc28955, nc28956, nc28957, nc28958, nc28959, nc28960, nc28961, nc28962, nc28963, nc28964, nc28965, nc28966, nc28967, nc28968, nc28969, nc28970, nc28971, nc28972, nc28973, nc28974, nc28975, nc28976, nc28977, nc28978, nc28979, nc28980, dw[46]}),
		.dipa (),
		.dipb (),
		.cea (net_719),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u372 (
		.sel (addra_pipe_0_net),
		.i0 (net_717),
		.i1 (net_721),
		.o (net_723)
	);
fifo2ram_emb_v1_AND u373 (
		.i0 (net_725),
		.i1 (net_724),
		.o (net_715)
	);
fifo2ram_emb_v1_AND u374 (
		.i0 (net_725),
		.i1 (ar[0]),
		.o (net_719)
	);
fifo2ram_emb_v1_NOT u375 (
		.i (ar[0]),
		.o (net_724)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_408 (
		.doa ({nc28981, nc28982, nc28983, nc28984, nc28985, nc28986, nc28987, nc28988, nc28989, nc28990, nc28991, nc28992, nc28993, nc28994, nc28995, nc28996, nc28997, nc28998, nc28999, nc29000, nc29001, nc29002, nc29003, nc29004, nc29005, nc29006, nc29007, nc29008, nc29009, nc29010, nc29011, nc29012, nc29013, nc29014, nc29015, nc29016, nc29017, nc29018, nc29019, nc29020, nc29021, nc29022, nc29023, nc29024, nc29025, nc29026, nc29027, nc29028, nc29029, nc29030, nc29031, nc29032, nc29033, nc29034, nc29035, nc29036, nc29037, nc29038, nc29039, nc29040, nc29041, nc29042, nc29043, net_728}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29044, nc29045, nc29046, nc29047, nc29048, nc29049, nc29050, nc29051, nc29052, nc29053, nc29054, nc29055, nc29056, nc29057, nc29058, nc29059, nc29060, nc29061, nc29062, nc29063, nc29064, nc29065, nc29066, nc29067, nc29068, nc29069, nc29070, nc29071, nc29072, nc29073, nc29074, nc29075, nc29076, nc29077, nc29078, nc29079, nc29080, nc29081, nc29082, nc29083, nc29084, nc29085, nc29086, nc29087, nc29088, nc29089, nc29090, nc29091, nc29092, nc29093, nc29094, nc29095, nc29096, nc29097, nc29098, nc29099, nc29100, nc29101, nc29102, nc29103, nc29104, nc29105, nc29106, dw[54]}),
		.dipa (),
		.dipb (),
		.cea (net_726),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_412 (
		.doa ({nc29107, nc29108, nc29109, nc29110, nc29111, nc29112, nc29113, nc29114, nc29115, nc29116, nc29117, nc29118, nc29119, nc29120, nc29121, nc29122, nc29123, nc29124, nc29125, nc29126, nc29127, nc29128, nc29129, nc29130, nc29131, nc29132, nc29133, nc29134, nc29135, nc29136, nc29137, nc29138, nc29139, nc29140, nc29141, nc29142, nc29143, nc29144, nc29145, nc29146, nc29147, nc29148, nc29149, nc29150, nc29151, nc29152, nc29153, nc29154, nc29155, nc29156, nc29157, nc29158, nc29159, nc29160, nc29161, nc29162, nc29163, nc29164, nc29165, nc29166, nc29167, nc29168, nc29169, net_732}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29170, nc29171, nc29172, nc29173, nc29174, nc29175, nc29176, nc29177, nc29178, nc29179, nc29180, nc29181, nc29182, nc29183, nc29184, nc29185, nc29186, nc29187, nc29188, nc29189, nc29190, nc29191, nc29192, nc29193, nc29194, nc29195, nc29196, nc29197, nc29198, nc29199, nc29200, nc29201, nc29202, nc29203, nc29204, nc29205, nc29206, nc29207, nc29208, nc29209, nc29210, nc29211, nc29212, nc29213, nc29214, nc29215, nc29216, nc29217, nc29218, nc29219, nc29220, nc29221, nc29222, nc29223, nc29224, nc29225, nc29226, nc29227, nc29228, nc29229, nc29230, nc29231, nc29232, dw[62]}),
		.dipa (),
		.dipb (),
		.cea (net_730),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u376 (
		.sel (addra_pipe_0_net),
		.i0 (net_728),
		.i1 (net_732),
		.o (net_734)
	);
fifo2ram_emb_v1_AND u377 (
		.i0 (net_736),
		.i1 (net_735),
		.o (net_726)
	);
fifo2ram_emb_v1_AND u378 (
		.i0 (net_736),
		.i1 (ar[0]),
		.o (net_730)
	);
fifo2ram_emb_v1_NOT u379 (
		.i (ar[0]),
		.o (net_735)
	);
fifo2ram_emb_v1_MUX u380 (
		.sel (addra_pipe_1_net),
		.i0 (net_723),
		.i1 (net_734),
		.o (net_737)
	);
fifo2ram_emb_v1_AND u381 (
		.i0 (net_739),
		.i1 (net_738),
		.o (net_725)
	);
fifo2ram_emb_v1_AND u382 (
		.i0 (net_739),
		.i1 (ar[1]),
		.o (net_736)
	);
fifo2ram_emb_v1_NOT u383 (
		.i (ar[1]),
		.o (net_738)
	);
fifo2ram_emb_v1_MUX u384 (
		.sel (addra_pipe_2_net),
		.i0 (net_712),
		.i1 (net_737),
		.o (net_740)
	);
fifo2ram_emb_v1_AND u385 (
		.i0 (net_742),
		.i1 (net_741),
		.o (net_714)
	);
fifo2ram_emb_v1_AND u386 (
		.i0 (net_742),
		.i1 (ar[2]),
		.o (net_739)
	);
fifo2ram_emb_v1_NOT u387 (
		.i (ar[2]),
		.o (net_741)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_416 (
		.doa ({nc29233, nc29234, nc29235, nc29236, nc29237, nc29238, nc29239, nc29240, nc29241, nc29242, nc29243, nc29244, nc29245, nc29246, nc29247, nc29248, nc29249, nc29250, nc29251, nc29252, nc29253, nc29254, nc29255, nc29256, nc29257, nc29258, nc29259, nc29260, nc29261, nc29262, nc29263, nc29264, nc29265, nc29266, nc29267, nc29268, nc29269, nc29270, nc29271, nc29272, nc29273, nc29274, nc29275, nc29276, nc29277, nc29278, nc29279, nc29280, nc29281, nc29282, nc29283, nc29284, nc29285, nc29286, nc29287, nc29288, nc29289, nc29290, nc29291, nc29292, nc29293, nc29294, nc29295, net_745}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29296, nc29297, nc29298, nc29299, nc29300, nc29301, nc29302, nc29303, nc29304, nc29305, nc29306, nc29307, nc29308, nc29309, nc29310, nc29311, nc29312, nc29313, nc29314, nc29315, nc29316, nc29317, nc29318, nc29319, nc29320, nc29321, nc29322, nc29323, nc29324, nc29325, nc29326, nc29327, nc29328, nc29329, nc29330, nc29331, nc29332, nc29333, nc29334, nc29335, nc29336, nc29337, nc29338, nc29339, nc29340, nc29341, nc29342, nc29343, nc29344, nc29345, nc29346, nc29347, nc29348, nc29349, nc29350, nc29351, nc29352, nc29353, nc29354, nc29355, nc29356, nc29357, nc29358, dw[70]}),
		.dipa (),
		.dipb (),
		.cea (net_743),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_420 (
		.doa ({nc29359, nc29360, nc29361, nc29362, nc29363, nc29364, nc29365, nc29366, nc29367, nc29368, nc29369, nc29370, nc29371, nc29372, nc29373, nc29374, nc29375, nc29376, nc29377, nc29378, nc29379, nc29380, nc29381, nc29382, nc29383, nc29384, nc29385, nc29386, nc29387, nc29388, nc29389, nc29390, nc29391, nc29392, nc29393, nc29394, nc29395, nc29396, nc29397, nc29398, nc29399, nc29400, nc29401, nc29402, nc29403, nc29404, nc29405, nc29406, nc29407, nc29408, nc29409, nc29410, nc29411, nc29412, nc29413, nc29414, nc29415, nc29416, nc29417, nc29418, nc29419, nc29420, nc29421, net_749}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29422, nc29423, nc29424, nc29425, nc29426, nc29427, nc29428, nc29429, nc29430, nc29431, nc29432, nc29433, nc29434, nc29435, nc29436, nc29437, nc29438, nc29439, nc29440, nc29441, nc29442, nc29443, nc29444, nc29445, nc29446, nc29447, nc29448, nc29449, nc29450, nc29451, nc29452, nc29453, nc29454, nc29455, nc29456, nc29457, nc29458, nc29459, nc29460, nc29461, nc29462, nc29463, nc29464, nc29465, nc29466, nc29467, nc29468, nc29469, nc29470, nc29471, nc29472, nc29473, nc29474, nc29475, nc29476, nc29477, nc29478, nc29479, nc29480, nc29481, nc29482, nc29483, nc29484, dw[78]}),
		.dipa (),
		.dipb (),
		.cea (net_747),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u388 (
		.sel (addra_pipe_0_net),
		.i0 (net_745),
		.i1 (net_749),
		.o (net_751)
	);
fifo2ram_emb_v1_AND u389 (
		.i0 (net_753),
		.i1 (net_752),
		.o (net_743)
	);
fifo2ram_emb_v1_AND u390 (
		.i0 (net_753),
		.i1 (ar[0]),
		.o (net_747)
	);
fifo2ram_emb_v1_NOT u391 (
		.i (ar[0]),
		.o (net_752)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_424 (
		.doa ({nc29485, nc29486, nc29487, nc29488, nc29489, nc29490, nc29491, nc29492, nc29493, nc29494, nc29495, nc29496, nc29497, nc29498, nc29499, nc29500, nc29501, nc29502, nc29503, nc29504, nc29505, nc29506, nc29507, nc29508, nc29509, nc29510, nc29511, nc29512, nc29513, nc29514, nc29515, nc29516, nc29517, nc29518, nc29519, nc29520, nc29521, nc29522, nc29523, nc29524, nc29525, nc29526, nc29527, nc29528, nc29529, nc29530, nc29531, nc29532, nc29533, nc29534, nc29535, nc29536, nc29537, nc29538, nc29539, nc29540, nc29541, nc29542, nc29543, nc29544, nc29545, nc29546, nc29547, net_756}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29548, nc29549, nc29550, nc29551, nc29552, nc29553, nc29554, nc29555, nc29556, nc29557, nc29558, nc29559, nc29560, nc29561, nc29562, nc29563, nc29564, nc29565, nc29566, nc29567, nc29568, nc29569, nc29570, nc29571, nc29572, nc29573, nc29574, nc29575, nc29576, nc29577, nc29578, nc29579, nc29580, nc29581, nc29582, nc29583, nc29584, nc29585, nc29586, nc29587, nc29588, nc29589, nc29590, nc29591, nc29592, nc29593, nc29594, nc29595, nc29596, nc29597, nc29598, nc29599, nc29600, nc29601, nc29602, nc29603, nc29604, nc29605, nc29606, nc29607, nc29608, nc29609, nc29610, dw[86]}),
		.dipa (),
		.dipb (),
		.cea (net_754),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_428 (
		.doa ({nc29611, nc29612, nc29613, nc29614, nc29615, nc29616, nc29617, nc29618, nc29619, nc29620, nc29621, nc29622, nc29623, nc29624, nc29625, nc29626, nc29627, nc29628, nc29629, nc29630, nc29631, nc29632, nc29633, nc29634, nc29635, nc29636, nc29637, nc29638, nc29639, nc29640, nc29641, nc29642, nc29643, nc29644, nc29645, nc29646, nc29647, nc29648, nc29649, nc29650, nc29651, nc29652, nc29653, nc29654, nc29655, nc29656, nc29657, nc29658, nc29659, nc29660, nc29661, nc29662, nc29663, nc29664, nc29665, nc29666, nc29667, nc29668, nc29669, nc29670, nc29671, nc29672, nc29673, net_760}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29674, nc29675, nc29676, nc29677, nc29678, nc29679, nc29680, nc29681, nc29682, nc29683, nc29684, nc29685, nc29686, nc29687, nc29688, nc29689, nc29690, nc29691, nc29692, nc29693, nc29694, nc29695, nc29696, nc29697, nc29698, nc29699, nc29700, nc29701, nc29702, nc29703, nc29704, nc29705, nc29706, nc29707, nc29708, nc29709, nc29710, nc29711, nc29712, nc29713, nc29714, nc29715, nc29716, nc29717, nc29718, nc29719, nc29720, nc29721, nc29722, nc29723, nc29724, nc29725, nc29726, nc29727, nc29728, nc29729, nc29730, nc29731, nc29732, nc29733, nc29734, nc29735, nc29736, dw[94]}),
		.dipa (),
		.dipb (),
		.cea (net_758),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u392 (
		.sel (addra_pipe_0_net),
		.i0 (net_756),
		.i1 (net_760),
		.o (net_762)
	);
fifo2ram_emb_v1_AND u393 (
		.i0 (net_764),
		.i1 (net_763),
		.o (net_754)
	);
fifo2ram_emb_v1_AND u394 (
		.i0 (net_764),
		.i1 (ar[0]),
		.o (net_758)
	);
fifo2ram_emb_v1_NOT u395 (
		.i (ar[0]),
		.o (net_763)
	);
fifo2ram_emb_v1_MUX u396 (
		.sel (addra_pipe_1_net),
		.i0 (net_751),
		.i1 (net_762),
		.o (net_765)
	);
fifo2ram_emb_v1_AND u397 (
		.i0 (net_767),
		.i1 (net_766),
		.o (net_753)
	);
fifo2ram_emb_v1_AND u398 (
		.i0 (net_767),
		.i1 (ar[1]),
		.o (net_764)
	);
fifo2ram_emb_v1_NOT u399 (
		.i (ar[1]),
		.o (net_766)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_432 (
		.doa ({nc29737, nc29738, nc29739, nc29740, nc29741, nc29742, nc29743, nc29744, nc29745, nc29746, nc29747, nc29748, nc29749, nc29750, nc29751, nc29752, nc29753, nc29754, nc29755, nc29756, nc29757, nc29758, nc29759, nc29760, nc29761, nc29762, nc29763, nc29764, nc29765, nc29766, nc29767, nc29768, nc29769, nc29770, nc29771, nc29772, nc29773, nc29774, nc29775, nc29776, nc29777, nc29778, nc29779, nc29780, nc29781, nc29782, nc29783, nc29784, nc29785, nc29786, nc29787, nc29788, nc29789, nc29790, nc29791, nc29792, nc29793, nc29794, nc29795, nc29796, nc29797, nc29798, nc29799, net_770}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29800, nc29801, nc29802, nc29803, nc29804, nc29805, nc29806, nc29807, nc29808, nc29809, nc29810, nc29811, nc29812, nc29813, nc29814, nc29815, nc29816, nc29817, nc29818, nc29819, nc29820, nc29821, nc29822, nc29823, nc29824, nc29825, nc29826, nc29827, nc29828, nc29829, nc29830, nc29831, nc29832, nc29833, nc29834, nc29835, nc29836, nc29837, nc29838, nc29839, nc29840, nc29841, nc29842, nc29843, nc29844, nc29845, nc29846, nc29847, nc29848, nc29849, nc29850, nc29851, nc29852, nc29853, nc29854, nc29855, nc29856, nc29857, nc29858, nc29859, nc29860, nc29861, nc29862, dw[102]}),
		.dipa (),
		.dipb (),
		.cea (net_768),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_436 (
		.doa ({nc29863, nc29864, nc29865, nc29866, nc29867, nc29868, nc29869, nc29870, nc29871, nc29872, nc29873, nc29874, nc29875, nc29876, nc29877, nc29878, nc29879, nc29880, nc29881, nc29882, nc29883, nc29884, nc29885, nc29886, nc29887, nc29888, nc29889, nc29890, nc29891, nc29892, nc29893, nc29894, nc29895, nc29896, nc29897, nc29898, nc29899, nc29900, nc29901, nc29902, nc29903, nc29904, nc29905, nc29906, nc29907, nc29908, nc29909, nc29910, nc29911, nc29912, nc29913, nc29914, nc29915, nc29916, nc29917, nc29918, nc29919, nc29920, nc29921, nc29922, nc29923, nc29924, nc29925, net_774}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc29926, nc29927, nc29928, nc29929, nc29930, nc29931, nc29932, nc29933, nc29934, nc29935, nc29936, nc29937, nc29938, nc29939, nc29940, nc29941, nc29942, nc29943, nc29944, nc29945, nc29946, nc29947, nc29948, nc29949, nc29950, nc29951, nc29952, nc29953, nc29954, nc29955, nc29956, nc29957, nc29958, nc29959, nc29960, nc29961, nc29962, nc29963, nc29964, nc29965, nc29966, nc29967, nc29968, nc29969, nc29970, nc29971, nc29972, nc29973, nc29974, nc29975, nc29976, nc29977, nc29978, nc29979, nc29980, nc29981, nc29982, nc29983, nc29984, nc29985, nc29986, nc29987, nc29988, dw[110]}),
		.dipa (),
		.dipb (),
		.cea (net_772),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u400 (
		.sel (addra_pipe_0_net),
		.i0 (net_770),
		.i1 (net_774),
		.o (net_776)
	);
fifo2ram_emb_v1_AND u401 (
		.i0 (net_778),
		.i1 (net_777),
		.o (net_768)
	);
fifo2ram_emb_v1_AND u402 (
		.i0 (net_778),
		.i1 (ar[0]),
		.o (net_772)
	);
fifo2ram_emb_v1_NOT u403 (
		.i (ar[0]),
		.o (net_777)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_440 (
		.doa ({nc29989, nc29990, nc29991, nc29992, nc29993, nc29994, nc29995, nc29996, nc29997, nc29998, nc29999, nc30000, nc30001, nc30002, nc30003, nc30004, nc30005, nc30006, nc30007, nc30008, nc30009, nc30010, nc30011, nc30012, nc30013, nc30014, nc30015, nc30016, nc30017, nc30018, nc30019, nc30020, nc30021, nc30022, nc30023, nc30024, nc30025, nc30026, nc30027, nc30028, nc30029, nc30030, nc30031, nc30032, nc30033, nc30034, nc30035, nc30036, nc30037, nc30038, nc30039, nc30040, nc30041, nc30042, nc30043, nc30044, nc30045, nc30046, nc30047, nc30048, nc30049, nc30050, nc30051, net_781}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30052, nc30053, nc30054, nc30055, nc30056, nc30057, nc30058, nc30059, nc30060, nc30061, nc30062, nc30063, nc30064, nc30065, nc30066, nc30067, nc30068, nc30069, nc30070, nc30071, nc30072, nc30073, nc30074, nc30075, nc30076, nc30077, nc30078, nc30079, nc30080, nc30081, nc30082, nc30083, nc30084, nc30085, nc30086, nc30087, nc30088, nc30089, nc30090, nc30091, nc30092, nc30093, nc30094, nc30095, nc30096, nc30097, nc30098, nc30099, nc30100, nc30101, nc30102, nc30103, nc30104, nc30105, nc30106, nc30107, nc30108, nc30109, nc30110, nc30111, nc30112, nc30113, nc30114, dw[118]}),
		.dipa (),
		.dipb (),
		.cea (net_779),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_444 (
		.doa ({nc30115, nc30116, nc30117, nc30118, nc30119, nc30120, nc30121, nc30122, nc30123, nc30124, nc30125, nc30126, nc30127, nc30128, nc30129, nc30130, nc30131, nc30132, nc30133, nc30134, nc30135, nc30136, nc30137, nc30138, nc30139, nc30140, nc30141, nc30142, nc30143, nc30144, nc30145, nc30146, nc30147, nc30148, nc30149, nc30150, nc30151, nc30152, nc30153, nc30154, nc30155, nc30156, nc30157, nc30158, nc30159, nc30160, nc30161, nc30162, nc30163, nc30164, nc30165, nc30166, nc30167, nc30168, nc30169, nc30170, nc30171, nc30172, nc30173, nc30174, nc30175, nc30176, nc30177, net_785}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30178, nc30179, nc30180, nc30181, nc30182, nc30183, nc30184, nc30185, nc30186, nc30187, nc30188, nc30189, nc30190, nc30191, nc30192, nc30193, nc30194, nc30195, nc30196, nc30197, nc30198, nc30199, nc30200, nc30201, nc30202, nc30203, nc30204, nc30205, nc30206, nc30207, nc30208, nc30209, nc30210, nc30211, nc30212, nc30213, nc30214, nc30215, nc30216, nc30217, nc30218, nc30219, nc30220, nc30221, nc30222, nc30223, nc30224, nc30225, nc30226, nc30227, nc30228, nc30229, nc30230, nc30231, nc30232, nc30233, nc30234, nc30235, nc30236, nc30237, nc30238, nc30239, nc30240, dw[126]}),
		.dipa (),
		.dipb (),
		.cea (net_783),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u404 (
		.sel (addra_pipe_0_net),
		.i0 (net_781),
		.i1 (net_785),
		.o (net_787)
	);
fifo2ram_emb_v1_AND u405 (
		.i0 (net_789),
		.i1 (net_788),
		.o (net_779)
	);
fifo2ram_emb_v1_AND u406 (
		.i0 (net_789),
		.i1 (ar[0]),
		.o (net_783)
	);
fifo2ram_emb_v1_NOT u407 (
		.i (ar[0]),
		.o (net_788)
	);
fifo2ram_emb_v1_MUX u408 (
		.sel (addra_pipe_1_net),
		.i0 (net_776),
		.i1 (net_787),
		.o (net_790)
	);
fifo2ram_emb_v1_AND u409 (
		.i0 (net_792),
		.i1 (net_791),
		.o (net_778)
	);
fifo2ram_emb_v1_AND u410 (
		.i0 (net_792),
		.i1 (ar[1]),
		.o (net_789)
	);
fifo2ram_emb_v1_NOT u411 (
		.i (ar[1]),
		.o (net_791)
	);
fifo2ram_emb_v1_MUX u412 (
		.sel (addra_pipe_2_net),
		.i0 (net_765),
		.i1 (net_790),
		.o (net_793)
	);
fifo2ram_emb_v1_AND u413 (
		.i0 (net_795),
		.i1 (net_794),
		.o (net_767)
	);
fifo2ram_emb_v1_AND u414 (
		.i0 (net_795),
		.i1 (ar[2]),
		.o (net_792)
	);
fifo2ram_emb_v1_NOT u415 (
		.i (ar[2]),
		.o (net_794)
	);
fifo2ram_emb_v1_MUX u416 (
		.sel (addra_pipe_3_net),
		.i0 (net_740),
		.i1 (net_793),
		.o (qr[6])
	);
fifo2ram_emb_v1_AND u417 (
		.i0 (cer),
		.i1 (net_797),
		.o (net_742)
	);
fifo2ram_emb_v1_AND u418 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_795)
	);
fifo2ram_emb_v1_NOT u419 (
		.i (ar[3]),
		.o (net_797)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_448 (
		.doa ({nc30241, nc30242, nc30243, nc30244, nc30245, nc30246, nc30247, nc30248, nc30249, nc30250, nc30251, nc30252, nc30253, nc30254, nc30255, nc30256, nc30257, nc30258, nc30259, nc30260, nc30261, nc30262, nc30263, nc30264, nc30265, nc30266, nc30267, nc30268, nc30269, nc30270, nc30271, nc30272, nc30273, nc30274, nc30275, nc30276, nc30277, nc30278, nc30279, nc30280, nc30281, nc30282, nc30283, nc30284, nc30285, nc30286, nc30287, nc30288, nc30289, nc30290, nc30291, nc30292, nc30293, nc30294, nc30295, nc30296, nc30297, nc30298, nc30299, nc30300, nc30301, nc30302, nc30303, net_801}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30304, nc30305, nc30306, nc30307, nc30308, nc30309, nc30310, nc30311, nc30312, nc30313, nc30314, nc30315, nc30316, nc30317, nc30318, nc30319, nc30320, nc30321, nc30322, nc30323, nc30324, nc30325, nc30326, nc30327, nc30328, nc30329, nc30330, nc30331, nc30332, nc30333, nc30334, nc30335, nc30336, nc30337, nc30338, nc30339, nc30340, nc30341, nc30342, nc30343, nc30344, nc30345, nc30346, nc30347, nc30348, nc30349, nc30350, nc30351, nc30352, nc30353, nc30354, nc30355, nc30356, nc30357, nc30358, nc30359, nc30360, nc30361, nc30362, nc30363, nc30364, nc30365, nc30366, dw[7]}),
		.dipa (),
		.dipb (),
		.cea (net_799),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_452 (
		.doa ({nc30367, nc30368, nc30369, nc30370, nc30371, nc30372, nc30373, nc30374, nc30375, nc30376, nc30377, nc30378, nc30379, nc30380, nc30381, nc30382, nc30383, nc30384, nc30385, nc30386, nc30387, nc30388, nc30389, nc30390, nc30391, nc30392, nc30393, nc30394, nc30395, nc30396, nc30397, nc30398, nc30399, nc30400, nc30401, nc30402, nc30403, nc30404, nc30405, nc30406, nc30407, nc30408, nc30409, nc30410, nc30411, nc30412, nc30413, nc30414, nc30415, nc30416, nc30417, nc30418, nc30419, nc30420, nc30421, nc30422, nc30423, nc30424, nc30425, nc30426, nc30427, nc30428, nc30429, net_805}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30430, nc30431, nc30432, nc30433, nc30434, nc30435, nc30436, nc30437, nc30438, nc30439, nc30440, nc30441, nc30442, nc30443, nc30444, nc30445, nc30446, nc30447, nc30448, nc30449, nc30450, nc30451, nc30452, nc30453, nc30454, nc30455, nc30456, nc30457, nc30458, nc30459, nc30460, nc30461, nc30462, nc30463, nc30464, nc30465, nc30466, nc30467, nc30468, nc30469, nc30470, nc30471, nc30472, nc30473, nc30474, nc30475, nc30476, nc30477, nc30478, nc30479, nc30480, nc30481, nc30482, nc30483, nc30484, nc30485, nc30486, nc30487, nc30488, nc30489, nc30490, nc30491, nc30492, dw[15]}),
		.dipa (),
		.dipb (),
		.cea (net_803),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u420 (
		.sel (addra_pipe_0_net),
		.i0 (net_801),
		.i1 (net_805),
		.o (net_807)
	);
fifo2ram_emb_v1_AND u421 (
		.i0 (net_809),
		.i1 (net_808),
		.o (net_799)
	);
fifo2ram_emb_v1_AND u422 (
		.i0 (net_809),
		.i1 (ar[0]),
		.o (net_803)
	);
fifo2ram_emb_v1_NOT u423 (
		.i (ar[0]),
		.o (net_808)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_456 (
		.doa ({nc30493, nc30494, nc30495, nc30496, nc30497, nc30498, nc30499, nc30500, nc30501, nc30502, nc30503, nc30504, nc30505, nc30506, nc30507, nc30508, nc30509, nc30510, nc30511, nc30512, nc30513, nc30514, nc30515, nc30516, nc30517, nc30518, nc30519, nc30520, nc30521, nc30522, nc30523, nc30524, nc30525, nc30526, nc30527, nc30528, nc30529, nc30530, nc30531, nc30532, nc30533, nc30534, nc30535, nc30536, nc30537, nc30538, nc30539, nc30540, nc30541, nc30542, nc30543, nc30544, nc30545, nc30546, nc30547, nc30548, nc30549, nc30550, nc30551, nc30552, nc30553, nc30554, nc30555, net_812}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30556, nc30557, nc30558, nc30559, nc30560, nc30561, nc30562, nc30563, nc30564, nc30565, nc30566, nc30567, nc30568, nc30569, nc30570, nc30571, nc30572, nc30573, nc30574, nc30575, nc30576, nc30577, nc30578, nc30579, nc30580, nc30581, nc30582, nc30583, nc30584, nc30585, nc30586, nc30587, nc30588, nc30589, nc30590, nc30591, nc30592, nc30593, nc30594, nc30595, nc30596, nc30597, nc30598, nc30599, nc30600, nc30601, nc30602, nc30603, nc30604, nc30605, nc30606, nc30607, nc30608, nc30609, nc30610, nc30611, nc30612, nc30613, nc30614, nc30615, nc30616, nc30617, nc30618, dw[23]}),
		.dipa (),
		.dipb (),
		.cea (net_810),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_460 (
		.doa ({nc30619, nc30620, nc30621, nc30622, nc30623, nc30624, nc30625, nc30626, nc30627, nc30628, nc30629, nc30630, nc30631, nc30632, nc30633, nc30634, nc30635, nc30636, nc30637, nc30638, nc30639, nc30640, nc30641, nc30642, nc30643, nc30644, nc30645, nc30646, nc30647, nc30648, nc30649, nc30650, nc30651, nc30652, nc30653, nc30654, nc30655, nc30656, nc30657, nc30658, nc30659, nc30660, nc30661, nc30662, nc30663, nc30664, nc30665, nc30666, nc30667, nc30668, nc30669, nc30670, nc30671, nc30672, nc30673, nc30674, nc30675, nc30676, nc30677, nc30678, nc30679, nc30680, nc30681, net_816}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30682, nc30683, nc30684, nc30685, nc30686, nc30687, nc30688, nc30689, nc30690, nc30691, nc30692, nc30693, nc30694, nc30695, nc30696, nc30697, nc30698, nc30699, nc30700, nc30701, nc30702, nc30703, nc30704, nc30705, nc30706, nc30707, nc30708, nc30709, nc30710, nc30711, nc30712, nc30713, nc30714, nc30715, nc30716, nc30717, nc30718, nc30719, nc30720, nc30721, nc30722, nc30723, nc30724, nc30725, nc30726, nc30727, nc30728, nc30729, nc30730, nc30731, nc30732, nc30733, nc30734, nc30735, nc30736, nc30737, nc30738, nc30739, nc30740, nc30741, nc30742, nc30743, nc30744, dw[31]}),
		.dipa (),
		.dipb (),
		.cea (net_814),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u424 (
		.sel (addra_pipe_0_net),
		.i0 (net_812),
		.i1 (net_816),
		.o (net_818)
	);
fifo2ram_emb_v1_AND u425 (
		.i0 (net_820),
		.i1 (net_819),
		.o (net_810)
	);
fifo2ram_emb_v1_AND u426 (
		.i0 (net_820),
		.i1 (ar[0]),
		.o (net_814)
	);
fifo2ram_emb_v1_NOT u427 (
		.i (ar[0]),
		.o (net_819)
	);
fifo2ram_emb_v1_MUX u428 (
		.sel (addra_pipe_1_net),
		.i0 (net_807),
		.i1 (net_818),
		.o (net_821)
	);
fifo2ram_emb_v1_AND u429 (
		.i0 (net_823),
		.i1 (net_822),
		.o (net_809)
	);
fifo2ram_emb_v1_AND u430 (
		.i0 (net_823),
		.i1 (ar[1]),
		.o (net_820)
	);
fifo2ram_emb_v1_NOT u431 (
		.i (ar[1]),
		.o (net_822)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_464 (
		.doa ({nc30745, nc30746, nc30747, nc30748, nc30749, nc30750, nc30751, nc30752, nc30753, nc30754, nc30755, nc30756, nc30757, nc30758, nc30759, nc30760, nc30761, nc30762, nc30763, nc30764, nc30765, nc30766, nc30767, nc30768, nc30769, nc30770, nc30771, nc30772, nc30773, nc30774, nc30775, nc30776, nc30777, nc30778, nc30779, nc30780, nc30781, nc30782, nc30783, nc30784, nc30785, nc30786, nc30787, nc30788, nc30789, nc30790, nc30791, nc30792, nc30793, nc30794, nc30795, nc30796, nc30797, nc30798, nc30799, nc30800, nc30801, nc30802, nc30803, nc30804, nc30805, nc30806, nc30807, net_826}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30808, nc30809, nc30810, nc30811, nc30812, nc30813, nc30814, nc30815, nc30816, nc30817, nc30818, nc30819, nc30820, nc30821, nc30822, nc30823, nc30824, nc30825, nc30826, nc30827, nc30828, nc30829, nc30830, nc30831, nc30832, nc30833, nc30834, nc30835, nc30836, nc30837, nc30838, nc30839, nc30840, nc30841, nc30842, nc30843, nc30844, nc30845, nc30846, nc30847, nc30848, nc30849, nc30850, nc30851, nc30852, nc30853, nc30854, nc30855, nc30856, nc30857, nc30858, nc30859, nc30860, nc30861, nc30862, nc30863, nc30864, nc30865, nc30866, nc30867, nc30868, nc30869, nc30870, dw[39]}),
		.dipa (),
		.dipb (),
		.cea (net_824),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_468 (
		.doa ({nc30871, nc30872, nc30873, nc30874, nc30875, nc30876, nc30877, nc30878, nc30879, nc30880, nc30881, nc30882, nc30883, nc30884, nc30885, nc30886, nc30887, nc30888, nc30889, nc30890, nc30891, nc30892, nc30893, nc30894, nc30895, nc30896, nc30897, nc30898, nc30899, nc30900, nc30901, nc30902, nc30903, nc30904, nc30905, nc30906, nc30907, nc30908, nc30909, nc30910, nc30911, nc30912, nc30913, nc30914, nc30915, nc30916, nc30917, nc30918, nc30919, nc30920, nc30921, nc30922, nc30923, nc30924, nc30925, nc30926, nc30927, nc30928, nc30929, nc30930, nc30931, nc30932, nc30933, net_830}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc30934, nc30935, nc30936, nc30937, nc30938, nc30939, nc30940, nc30941, nc30942, nc30943, nc30944, nc30945, nc30946, nc30947, nc30948, nc30949, nc30950, nc30951, nc30952, nc30953, nc30954, nc30955, nc30956, nc30957, nc30958, nc30959, nc30960, nc30961, nc30962, nc30963, nc30964, nc30965, nc30966, nc30967, nc30968, nc30969, nc30970, nc30971, nc30972, nc30973, nc30974, nc30975, nc30976, nc30977, nc30978, nc30979, nc30980, nc30981, nc30982, nc30983, nc30984, nc30985, nc30986, nc30987, nc30988, nc30989, nc30990, nc30991, nc30992, nc30993, nc30994, nc30995, nc30996, dw[47]}),
		.dipa (),
		.dipb (),
		.cea (net_828),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u432 (
		.sel (addra_pipe_0_net),
		.i0 (net_826),
		.i1 (net_830),
		.o (net_832)
	);
fifo2ram_emb_v1_AND u433 (
		.i0 (net_834),
		.i1 (net_833),
		.o (net_824)
	);
fifo2ram_emb_v1_AND u434 (
		.i0 (net_834),
		.i1 (ar[0]),
		.o (net_828)
	);
fifo2ram_emb_v1_NOT u435 (
		.i (ar[0]),
		.o (net_833)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_472 (
		.doa ({nc30997, nc30998, nc30999, nc31000, nc31001, nc31002, nc31003, nc31004, nc31005, nc31006, nc31007, nc31008, nc31009, nc31010, nc31011, nc31012, nc31013, nc31014, nc31015, nc31016, nc31017, nc31018, nc31019, nc31020, nc31021, nc31022, nc31023, nc31024, nc31025, nc31026, nc31027, nc31028, nc31029, nc31030, nc31031, nc31032, nc31033, nc31034, nc31035, nc31036, nc31037, nc31038, nc31039, nc31040, nc31041, nc31042, nc31043, nc31044, nc31045, nc31046, nc31047, nc31048, nc31049, nc31050, nc31051, nc31052, nc31053, nc31054, nc31055, nc31056, nc31057, nc31058, nc31059, net_837}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31060, nc31061, nc31062, nc31063, nc31064, nc31065, nc31066, nc31067, nc31068, nc31069, nc31070, nc31071, nc31072, nc31073, nc31074, nc31075, nc31076, nc31077, nc31078, nc31079, nc31080, nc31081, nc31082, nc31083, nc31084, nc31085, nc31086, nc31087, nc31088, nc31089, nc31090, nc31091, nc31092, nc31093, nc31094, nc31095, nc31096, nc31097, nc31098, nc31099, nc31100, nc31101, nc31102, nc31103, nc31104, nc31105, nc31106, nc31107, nc31108, nc31109, nc31110, nc31111, nc31112, nc31113, nc31114, nc31115, nc31116, nc31117, nc31118, nc31119, nc31120, nc31121, nc31122, dw[55]}),
		.dipa (),
		.dipb (),
		.cea (net_835),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_476 (
		.doa ({nc31123, nc31124, nc31125, nc31126, nc31127, nc31128, nc31129, nc31130, nc31131, nc31132, nc31133, nc31134, nc31135, nc31136, nc31137, nc31138, nc31139, nc31140, nc31141, nc31142, nc31143, nc31144, nc31145, nc31146, nc31147, nc31148, nc31149, nc31150, nc31151, nc31152, nc31153, nc31154, nc31155, nc31156, nc31157, nc31158, nc31159, nc31160, nc31161, nc31162, nc31163, nc31164, nc31165, nc31166, nc31167, nc31168, nc31169, nc31170, nc31171, nc31172, nc31173, nc31174, nc31175, nc31176, nc31177, nc31178, nc31179, nc31180, nc31181, nc31182, nc31183, nc31184, nc31185, net_841}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31186, nc31187, nc31188, nc31189, nc31190, nc31191, nc31192, nc31193, nc31194, nc31195, nc31196, nc31197, nc31198, nc31199, nc31200, nc31201, nc31202, nc31203, nc31204, nc31205, nc31206, nc31207, nc31208, nc31209, nc31210, nc31211, nc31212, nc31213, nc31214, nc31215, nc31216, nc31217, nc31218, nc31219, nc31220, nc31221, nc31222, nc31223, nc31224, nc31225, nc31226, nc31227, nc31228, nc31229, nc31230, nc31231, nc31232, nc31233, nc31234, nc31235, nc31236, nc31237, nc31238, nc31239, nc31240, nc31241, nc31242, nc31243, nc31244, nc31245, nc31246, nc31247, nc31248, dw[63]}),
		.dipa (),
		.dipb (),
		.cea (net_839),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u436 (
		.sel (addra_pipe_0_net),
		.i0 (net_837),
		.i1 (net_841),
		.o (net_843)
	);
fifo2ram_emb_v1_AND u437 (
		.i0 (net_845),
		.i1 (net_844),
		.o (net_835)
	);
fifo2ram_emb_v1_AND u438 (
		.i0 (net_845),
		.i1 (ar[0]),
		.o (net_839)
	);
fifo2ram_emb_v1_NOT u439 (
		.i (ar[0]),
		.o (net_844)
	);
fifo2ram_emb_v1_MUX u440 (
		.sel (addra_pipe_1_net),
		.i0 (net_832),
		.i1 (net_843),
		.o (net_846)
	);
fifo2ram_emb_v1_AND u441 (
		.i0 (net_848),
		.i1 (net_847),
		.o (net_834)
	);
fifo2ram_emb_v1_AND u442 (
		.i0 (net_848),
		.i1 (ar[1]),
		.o (net_845)
	);
fifo2ram_emb_v1_NOT u443 (
		.i (ar[1]),
		.o (net_847)
	);
fifo2ram_emb_v1_MUX u444 (
		.sel (addra_pipe_2_net),
		.i0 (net_821),
		.i1 (net_846),
		.o (net_849)
	);
fifo2ram_emb_v1_AND u445 (
		.i0 (net_851),
		.i1 (net_850),
		.o (net_823)
	);
fifo2ram_emb_v1_AND u446 (
		.i0 (net_851),
		.i1 (ar[2]),
		.o (net_848)
	);
fifo2ram_emb_v1_NOT u447 (
		.i (ar[2]),
		.o (net_850)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_480 (
		.doa ({nc31249, nc31250, nc31251, nc31252, nc31253, nc31254, nc31255, nc31256, nc31257, nc31258, nc31259, nc31260, nc31261, nc31262, nc31263, nc31264, nc31265, nc31266, nc31267, nc31268, nc31269, nc31270, nc31271, nc31272, nc31273, nc31274, nc31275, nc31276, nc31277, nc31278, nc31279, nc31280, nc31281, nc31282, nc31283, nc31284, nc31285, nc31286, nc31287, nc31288, nc31289, nc31290, nc31291, nc31292, nc31293, nc31294, nc31295, nc31296, nc31297, nc31298, nc31299, nc31300, nc31301, nc31302, nc31303, nc31304, nc31305, nc31306, nc31307, nc31308, nc31309, nc31310, nc31311, net_854}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31312, nc31313, nc31314, nc31315, nc31316, nc31317, nc31318, nc31319, nc31320, nc31321, nc31322, nc31323, nc31324, nc31325, nc31326, nc31327, nc31328, nc31329, nc31330, nc31331, nc31332, nc31333, nc31334, nc31335, nc31336, nc31337, nc31338, nc31339, nc31340, nc31341, nc31342, nc31343, nc31344, nc31345, nc31346, nc31347, nc31348, nc31349, nc31350, nc31351, nc31352, nc31353, nc31354, nc31355, nc31356, nc31357, nc31358, nc31359, nc31360, nc31361, nc31362, nc31363, nc31364, nc31365, nc31366, nc31367, nc31368, nc31369, nc31370, nc31371, nc31372, nc31373, nc31374, dw[71]}),
		.dipa (),
		.dipb (),
		.cea (net_852),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_484 (
		.doa ({nc31375, nc31376, nc31377, nc31378, nc31379, nc31380, nc31381, nc31382, nc31383, nc31384, nc31385, nc31386, nc31387, nc31388, nc31389, nc31390, nc31391, nc31392, nc31393, nc31394, nc31395, nc31396, nc31397, nc31398, nc31399, nc31400, nc31401, nc31402, nc31403, nc31404, nc31405, nc31406, nc31407, nc31408, nc31409, nc31410, nc31411, nc31412, nc31413, nc31414, nc31415, nc31416, nc31417, nc31418, nc31419, nc31420, nc31421, nc31422, nc31423, nc31424, nc31425, nc31426, nc31427, nc31428, nc31429, nc31430, nc31431, nc31432, nc31433, nc31434, nc31435, nc31436, nc31437, net_858}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31438, nc31439, nc31440, nc31441, nc31442, nc31443, nc31444, nc31445, nc31446, nc31447, nc31448, nc31449, nc31450, nc31451, nc31452, nc31453, nc31454, nc31455, nc31456, nc31457, nc31458, nc31459, nc31460, nc31461, nc31462, nc31463, nc31464, nc31465, nc31466, nc31467, nc31468, nc31469, nc31470, nc31471, nc31472, nc31473, nc31474, nc31475, nc31476, nc31477, nc31478, nc31479, nc31480, nc31481, nc31482, nc31483, nc31484, nc31485, nc31486, nc31487, nc31488, nc31489, nc31490, nc31491, nc31492, nc31493, nc31494, nc31495, nc31496, nc31497, nc31498, nc31499, nc31500, dw[79]}),
		.dipa (),
		.dipb (),
		.cea (net_856),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u448 (
		.sel (addra_pipe_0_net),
		.i0 (net_854),
		.i1 (net_858),
		.o (net_860)
	);
fifo2ram_emb_v1_AND u449 (
		.i0 (net_862),
		.i1 (net_861),
		.o (net_852)
	);
fifo2ram_emb_v1_AND u450 (
		.i0 (net_862),
		.i1 (ar[0]),
		.o (net_856)
	);
fifo2ram_emb_v1_NOT u451 (
		.i (ar[0]),
		.o (net_861)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_488 (
		.doa ({nc31501, nc31502, nc31503, nc31504, nc31505, nc31506, nc31507, nc31508, nc31509, nc31510, nc31511, nc31512, nc31513, nc31514, nc31515, nc31516, nc31517, nc31518, nc31519, nc31520, nc31521, nc31522, nc31523, nc31524, nc31525, nc31526, nc31527, nc31528, nc31529, nc31530, nc31531, nc31532, nc31533, nc31534, nc31535, nc31536, nc31537, nc31538, nc31539, nc31540, nc31541, nc31542, nc31543, nc31544, nc31545, nc31546, nc31547, nc31548, nc31549, nc31550, nc31551, nc31552, nc31553, nc31554, nc31555, nc31556, nc31557, nc31558, nc31559, nc31560, nc31561, nc31562, nc31563, net_865}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31564, nc31565, nc31566, nc31567, nc31568, nc31569, nc31570, nc31571, nc31572, nc31573, nc31574, nc31575, nc31576, nc31577, nc31578, nc31579, nc31580, nc31581, nc31582, nc31583, nc31584, nc31585, nc31586, nc31587, nc31588, nc31589, nc31590, nc31591, nc31592, nc31593, nc31594, nc31595, nc31596, nc31597, nc31598, nc31599, nc31600, nc31601, nc31602, nc31603, nc31604, nc31605, nc31606, nc31607, nc31608, nc31609, nc31610, nc31611, nc31612, nc31613, nc31614, nc31615, nc31616, nc31617, nc31618, nc31619, nc31620, nc31621, nc31622, nc31623, nc31624, nc31625, nc31626, dw[87]}),
		.dipa (),
		.dipb (),
		.cea (net_863),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_492 (
		.doa ({nc31627, nc31628, nc31629, nc31630, nc31631, nc31632, nc31633, nc31634, nc31635, nc31636, nc31637, nc31638, nc31639, nc31640, nc31641, nc31642, nc31643, nc31644, nc31645, nc31646, nc31647, nc31648, nc31649, nc31650, nc31651, nc31652, nc31653, nc31654, nc31655, nc31656, nc31657, nc31658, nc31659, nc31660, nc31661, nc31662, nc31663, nc31664, nc31665, nc31666, nc31667, nc31668, nc31669, nc31670, nc31671, nc31672, nc31673, nc31674, nc31675, nc31676, nc31677, nc31678, nc31679, nc31680, nc31681, nc31682, nc31683, nc31684, nc31685, nc31686, nc31687, nc31688, nc31689, net_869}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31690, nc31691, nc31692, nc31693, nc31694, nc31695, nc31696, nc31697, nc31698, nc31699, nc31700, nc31701, nc31702, nc31703, nc31704, nc31705, nc31706, nc31707, nc31708, nc31709, nc31710, nc31711, nc31712, nc31713, nc31714, nc31715, nc31716, nc31717, nc31718, nc31719, nc31720, nc31721, nc31722, nc31723, nc31724, nc31725, nc31726, nc31727, nc31728, nc31729, nc31730, nc31731, nc31732, nc31733, nc31734, nc31735, nc31736, nc31737, nc31738, nc31739, nc31740, nc31741, nc31742, nc31743, nc31744, nc31745, nc31746, nc31747, nc31748, nc31749, nc31750, nc31751, nc31752, dw[95]}),
		.dipa (),
		.dipb (),
		.cea (net_867),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u452 (
		.sel (addra_pipe_0_net),
		.i0 (net_865),
		.i1 (net_869),
		.o (net_871)
	);
fifo2ram_emb_v1_AND u453 (
		.i0 (net_873),
		.i1 (net_872),
		.o (net_863)
	);
fifo2ram_emb_v1_AND u454 (
		.i0 (net_873),
		.i1 (ar[0]),
		.o (net_867)
	);
fifo2ram_emb_v1_NOT u455 (
		.i (ar[0]),
		.o (net_872)
	);
fifo2ram_emb_v1_MUX u456 (
		.sel (addra_pipe_1_net),
		.i0 (net_860),
		.i1 (net_871),
		.o (net_874)
	);
fifo2ram_emb_v1_AND u457 (
		.i0 (net_876),
		.i1 (net_875),
		.o (net_862)
	);
fifo2ram_emb_v1_AND u458 (
		.i0 (net_876),
		.i1 (ar[1]),
		.o (net_873)
	);
fifo2ram_emb_v1_NOT u459 (
		.i (ar[1]),
		.o (net_875)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_496 (
		.doa ({nc31753, nc31754, nc31755, nc31756, nc31757, nc31758, nc31759, nc31760, nc31761, nc31762, nc31763, nc31764, nc31765, nc31766, nc31767, nc31768, nc31769, nc31770, nc31771, nc31772, nc31773, nc31774, nc31775, nc31776, nc31777, nc31778, nc31779, nc31780, nc31781, nc31782, nc31783, nc31784, nc31785, nc31786, nc31787, nc31788, nc31789, nc31790, nc31791, nc31792, nc31793, nc31794, nc31795, nc31796, nc31797, nc31798, nc31799, nc31800, nc31801, nc31802, nc31803, nc31804, nc31805, nc31806, nc31807, nc31808, nc31809, nc31810, nc31811, nc31812, nc31813, nc31814, nc31815, net_879}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31816, nc31817, nc31818, nc31819, nc31820, nc31821, nc31822, nc31823, nc31824, nc31825, nc31826, nc31827, nc31828, nc31829, nc31830, nc31831, nc31832, nc31833, nc31834, nc31835, nc31836, nc31837, nc31838, nc31839, nc31840, nc31841, nc31842, nc31843, nc31844, nc31845, nc31846, nc31847, nc31848, nc31849, nc31850, nc31851, nc31852, nc31853, nc31854, nc31855, nc31856, nc31857, nc31858, nc31859, nc31860, nc31861, nc31862, nc31863, nc31864, nc31865, nc31866, nc31867, nc31868, nc31869, nc31870, nc31871, nc31872, nc31873, nc31874, nc31875, nc31876, nc31877, nc31878, dw[103]}),
		.dipa (),
		.dipb (),
		.cea (net_877),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_500 (
		.doa ({nc31879, nc31880, nc31881, nc31882, nc31883, nc31884, nc31885, nc31886, nc31887, nc31888, nc31889, nc31890, nc31891, nc31892, nc31893, nc31894, nc31895, nc31896, nc31897, nc31898, nc31899, nc31900, nc31901, nc31902, nc31903, nc31904, nc31905, nc31906, nc31907, nc31908, nc31909, nc31910, nc31911, nc31912, nc31913, nc31914, nc31915, nc31916, nc31917, nc31918, nc31919, nc31920, nc31921, nc31922, nc31923, nc31924, nc31925, nc31926, nc31927, nc31928, nc31929, nc31930, nc31931, nc31932, nc31933, nc31934, nc31935, nc31936, nc31937, nc31938, nc31939, nc31940, nc31941, net_883}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc31942, nc31943, nc31944, nc31945, nc31946, nc31947, nc31948, nc31949, nc31950, nc31951, nc31952, nc31953, nc31954, nc31955, nc31956, nc31957, nc31958, nc31959, nc31960, nc31961, nc31962, nc31963, nc31964, nc31965, nc31966, nc31967, nc31968, nc31969, nc31970, nc31971, nc31972, nc31973, nc31974, nc31975, nc31976, nc31977, nc31978, nc31979, nc31980, nc31981, nc31982, nc31983, nc31984, nc31985, nc31986, nc31987, nc31988, nc31989, nc31990, nc31991, nc31992, nc31993, nc31994, nc31995, nc31996, nc31997, nc31998, nc31999, nc32000, nc32001, nc32002, nc32003, nc32004, dw[111]}),
		.dipa (),
		.dipb (),
		.cea (net_881),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u460 (
		.sel (addra_pipe_0_net),
		.i0 (net_879),
		.i1 (net_883),
		.o (net_885)
	);
fifo2ram_emb_v1_AND u461 (
		.i0 (net_887),
		.i1 (net_886),
		.o (net_877)
	);
fifo2ram_emb_v1_AND u462 (
		.i0 (net_887),
		.i1 (ar[0]),
		.o (net_881)
	);
fifo2ram_emb_v1_NOT u463 (
		.i (ar[0]),
		.o (net_886)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_504 (
		.doa ({nc32005, nc32006, nc32007, nc32008, nc32009, nc32010, nc32011, nc32012, nc32013, nc32014, nc32015, nc32016, nc32017, nc32018, nc32019, nc32020, nc32021, nc32022, nc32023, nc32024, nc32025, nc32026, nc32027, nc32028, nc32029, nc32030, nc32031, nc32032, nc32033, nc32034, nc32035, nc32036, nc32037, nc32038, nc32039, nc32040, nc32041, nc32042, nc32043, nc32044, nc32045, nc32046, nc32047, nc32048, nc32049, nc32050, nc32051, nc32052, nc32053, nc32054, nc32055, nc32056, nc32057, nc32058, nc32059, nc32060, nc32061, nc32062, nc32063, nc32064, nc32065, nc32066, nc32067, net_890}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc32068, nc32069, nc32070, nc32071, nc32072, nc32073, nc32074, nc32075, nc32076, nc32077, nc32078, nc32079, nc32080, nc32081, nc32082, nc32083, nc32084, nc32085, nc32086, nc32087, nc32088, nc32089, nc32090, nc32091, nc32092, nc32093, nc32094, nc32095, nc32096, nc32097, nc32098, nc32099, nc32100, nc32101, nc32102, nc32103, nc32104, nc32105, nc32106, nc32107, nc32108, nc32109, nc32110, nc32111, nc32112, nc32113, nc32114, nc32115, nc32116, nc32117, nc32118, nc32119, nc32120, nc32121, nc32122, nc32123, nc32124, nc32125, nc32126, nc32127, nc32128, nc32129, nc32130, dw[119]}),
		.dipa (),
		.dipb (),
		.cea (net_888),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
EMB18K #(
		.clka_inv (1'b0),
		.clkb_inv (1'b0),
		.eccreaden (1'b0),
		.eccwriteen (1'b0),
		.emb5k_1_init_file (""),
		.emb5k_2_init_file (""),
		.emb5k_3_init_file (""),
		.emb5k_4_init_file (""),
		.extension_mode ("power"),
		.init_file ("none"),
		.outreg_a (1'b0),
		.outreg_b (1'b0),
		.rammode ("sdp"),
		.use_parity (1'b0),
		.width_a (1),
		.width_b (1),
		.writemode_a ("write_first"),
		.writemode_b ("write_first")
	)
	emb_508 (
		.doa ({nc32131, nc32132, nc32133, nc32134, nc32135, nc32136, nc32137, nc32138, nc32139, nc32140, nc32141, nc32142, nc32143, nc32144, nc32145, nc32146, nc32147, nc32148, nc32149, nc32150, nc32151, nc32152, nc32153, nc32154, nc32155, nc32156, nc32157, nc32158, nc32159, nc32160, nc32161, nc32162, nc32163, nc32164, nc32165, nc32166, nc32167, nc32168, nc32169, nc32170, nc32171, nc32172, nc32173, nc32174, nc32175, nc32176, nc32177, nc32178, nc32179, nc32180, nc32181, nc32182, nc32183, nc32184, nc32185, nc32186, nc32187, nc32188, nc32189, nc32190, nc32191, nc32192, nc32193, net_894}),
		.dob (),
		.dopa (),
		.dopb (),
		.addra ({ar[17], ar[16], ar[15], ar[14], ar[13], ar[12], ar[11], ar[10], ar[9], ar[8], ar[7], ar[6], ar[5], ar[4]}),
		.addrb ({aw[13], aw[12], aw[11], aw[10], aw[9], aw[8], aw[7], aw[6], aw[5], aw[4], aw[3], aw[2], aw[1], aw[0]}),
		.clka (clkr),
		.clkb (clkw),
		.dia (),
		.dib ({nc32194, nc32195, nc32196, nc32197, nc32198, nc32199, nc32200, nc32201, nc32202, nc32203, nc32204, nc32205, nc32206, nc32207, nc32208, nc32209, nc32210, nc32211, nc32212, nc32213, nc32214, nc32215, nc32216, nc32217, nc32218, nc32219, nc32220, nc32221, nc32222, nc32223, nc32224, nc32225, nc32226, nc32227, nc32228, nc32229, nc32230, nc32231, nc32232, nc32233, nc32234, nc32235, nc32236, nc32237, nc32238, nc32239, nc32240, nc32241, nc32242, nc32243, nc32244, nc32245, nc32246, nc32247, nc32248, nc32249, nc32250, nc32251, nc32252, nc32253, nc32254, nc32255, nc32256, dw[127]}),
		.dipa (),
		.dipb (),
		.cea (net_892),
		.ceb (cew),
		.regcea (vcc_net),
		.regceb (),
		.regsra (rstnr),
		.regsrb (),
		.wea ({gnd_net, gnd_net, gnd_net, gnd_net}),
		.web ({vcc_net, vcc_net, vcc_net, vcc_net}),
		.eccoutdberr (),
		.eccoutsberr (),
		.eccreadaddr (),
		.eccindberr (gnd_net),
		.eccinsberr (gnd_net)
	);
fifo2ram_emb_v1_MUX u464 (
		.sel (addra_pipe_0_net),
		.i0 (net_890),
		.i1 (net_894),
		.o (net_896)
	);
fifo2ram_emb_v1_AND u465 (
		.i0 (net_898),
		.i1 (net_897),
		.o (net_888)
	);
fifo2ram_emb_v1_AND u466 (
		.i0 (net_898),
		.i1 (ar[0]),
		.o (net_892)
	);
fifo2ram_emb_v1_NOT u467 (
		.i (ar[0]),
		.o (net_897)
	);
fifo2ram_emb_v1_MUX u468 (
		.sel (addra_pipe_1_net),
		.i0 (net_885),
		.i1 (net_896),
		.o (net_899)
	);
fifo2ram_emb_v1_AND u469 (
		.i0 (net_901),
		.i1 (net_900),
		.o (net_887)
	);
fifo2ram_emb_v1_AND u470 (
		.i0 (net_901),
		.i1 (ar[1]),
		.o (net_898)
	);
fifo2ram_emb_v1_NOT u471 (
		.i (ar[1]),
		.o (net_900)
	);
fifo2ram_emb_v1_MUX u472 (
		.sel (addra_pipe_2_net),
		.i0 (net_874),
		.i1 (net_899),
		.o (net_902)
	);
fifo2ram_emb_v1_AND u473 (
		.i0 (net_904),
		.i1 (net_903),
		.o (net_876)
	);
fifo2ram_emb_v1_AND u474 (
		.i0 (net_904),
		.i1 (ar[2]),
		.o (net_901)
	);
fifo2ram_emb_v1_NOT u475 (
		.i (ar[2]),
		.o (net_903)
	);
fifo2ram_emb_v1_MUX u476 (
		.sel (addra_pipe_3_net),
		.i0 (net_849),
		.i1 (net_902),
		.o (qr[7])
	);
fifo2ram_emb_v1_AND u477 (
		.i0 (cer),
		.i1 (net_906),
		.o (net_851)
	);
fifo2ram_emb_v1_AND u478 (
		.i0 (cer),
		.i1 (ar[3]),
		.o (net_904)
	);
fifo2ram_emb_v1_NOT u479 (
		.i (ar[3]),
		.o (net_906)
	);

endmodule
module fifo2ram_emb_v1_ADDR_PIPE_A (clk, ena, i, o);
input clk;
input ena;
input i;
output o;



reg r0;
always @(posedge clk) begin
	if (ena) r0 <= i;
end
assign o = r0;

endmodule
module fifo2ram_emb_v1_MUX (sel, i0, i1, o);
input sel;
input i0;
input i1;
output o;



assign o = sel? i1 : i0;

endmodule
module fifo2ram_emb_v1_AND (i0, i1, o);
input i0;
input i1;
output o;



assign o = i0 & i1;

endmodule
module fifo2ram_emb_v1_NOT (i, o);
input i;
output o;



assign o = ~i;

endmodule
