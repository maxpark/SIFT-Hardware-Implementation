`timescale 1ns / 1ps


module local_gau_rom
(
    input   [7:0]       a,  // Addr.
	output  reg [7:0]	spo // Data.
);
	
	always @(*) begin
		case (a)
			000: spo = 8'h0;
            001: spo = 8'h1;
            002: spo = 8'h1;
            003: spo = 8'h1;
            004: spo = 8'h1;
            005: spo = 8'h2;
            006: spo = 8'h2;
            007: spo = 8'h2;
            008: spo = 8'h2;
            009: spo = 8'h2;
            010: spo = 8'h2;
            011: spo = 8'h1;
            012: spo = 8'h1;
            013: spo = 8'h1;
            014: spo = 8'h1;
            015: spo = 8'h0;
            016: spo = 8'h1;
            017: spo = 8'h1;
            018: spo = 8'h1;
            019: spo = 8'h2;
            020: spo = 8'h2;
            021: spo = 8'h2;
            022: spo = 8'h3;
            023: spo = 8'h3;
            024: spo = 8'h3;
            025: spo = 8'h3;
            026: spo = 8'h2;
            027: spo = 8'h2;
            028: spo = 8'h2;
            029: spo = 8'h1;
            030: spo = 8'h1;
            031: spo = 8'h1;
            032: spo = 8'h1;
            033: spo = 8'h1;
            034: spo = 8'h2;
            035: spo = 8'h2;
            036: spo = 8'h3;
            037: spo = 8'h4;
            038: spo = 8'h4;
            039: spo = 8'h4;
            040: spo = 8'h4;
            041: spo = 8'h4;
            042: spo = 8'h4;
            043: spo = 8'h3;
            044: spo = 8'h2;
            045: spo = 8'h2;
            046: spo = 8'h1;
            047: spo = 8'h1;
            048: spo = 8'h1;
            049: spo = 8'h2;
            050: spo = 8'h2;
            051: spo = 8'h3;
            052: spo = 8'h4;
            053: spo = 8'h5;
            054: spo = 8'h6;
            055: spo = 8'h6;
            056: spo = 8'h6;
            057: spo = 8'h6;
            058: spo = 8'h5;
            059: spo = 8'h4;
            060: spo = 8'h3;
            061: spo = 8'h2;
            062: spo = 8'h2;
            063: spo = 8'h1;
            064: spo = 8'h1;
            065: spo = 8'h2;
            066: spo = 8'h3;
            067: spo = 8'h4;
            068: spo = 8'h5;
            069: spo = 8'h6;
            070: spo = 8'h7;
            071: spo = 8'h8;
            072: spo = 8'h8;
            073: spo = 8'h7;
            074: spo = 8'h6;
            075: spo = 8'h5;
            076: spo = 8'h4;
            077: spo = 8'h3;
            078: spo = 8'h2;
            079: spo = 8'h1;
            080: spo = 8'h2;
            081: spo = 8'h2;
            082: spo = 8'h4;
            083: spo = 8'h5;
            084: spo = 8'h6;
            085: spo = 8'h8;
            086: spo = 8'h9;
            087: spo = 8'h9;
            088: spo = 8'h9;
            089: spo = 8'h9;
            090: spo = 8'h8;
            091: spo = 8'h6;
            092: spo = 8'h5;
            093: spo = 8'h4;
            094: spo = 8'h2;
            095: spo = 8'h2;
            096: spo = 8'h2;
            097: spo = 8'h3;
            098: spo = 8'h4;
            099: spo = 8'h6;
            100: spo = 8'h7;
            101: spo = 8'h9;
            102: spo = 8'ha;
            103: spo = 8'ha;
            104: spo = 8'ha;
            105: spo = 8'ha;
            106: spo = 8'h9;
            107: spo = 8'h7;
            108: spo = 8'h6;
            109: spo = 8'h4;
            110: spo = 8'h3;
            111: spo = 8'h2;
            112: spo = 8'h2;
            113: spo = 8'h3;
            114: spo = 8'h4;
            115: spo = 8'h6;
            116: spo = 8'h8;
            117: spo = 8'h9;
            118: spo = 8'ha;
            119: spo = 8'hb;
            120: spo = 8'hb;
            121: spo = 8'ha;
            122: spo = 8'h9;
            123: spo = 8'h8;
            124: spo = 8'h6;
            125: spo = 8'h4;
            126: spo = 8'h3;
            127: spo = 8'h2;
            128: spo = 8'h2;
            129: spo = 8'h3;
            130: spo = 8'h4;
            131: spo = 8'h6;
            132: spo = 8'h8;
            133: spo = 8'h9;
            134: spo = 8'ha;
            135: spo = 8'hb;
            136: spo = 8'hb;
            137: spo = 8'ha;
            138: spo = 8'h9;
            139: spo = 8'h8;
            140: spo = 8'h6;
            141: spo = 8'h4;
            142: spo = 8'h3;
            143: spo = 8'h2;
            144: spo = 8'h2;
            145: spo = 8'h3;
            146: spo = 8'h4;
            147: spo = 8'h6;
            148: spo = 8'h7;
            149: spo = 8'h9;
            150: spo = 8'ha;
            151: spo = 8'ha;
            152: spo = 8'ha;
            153: spo = 8'ha;
            154: spo = 8'h9;
            155: spo = 8'h7;
            156: spo = 8'h6;
            157: spo = 8'h4;
            158: spo = 8'h3;
            159: spo = 8'h2;
            160: spo = 8'h2;
            161: spo = 8'h2;
            162: spo = 8'h4;
            163: spo = 8'h5;
            164: spo = 8'h6;
            165: spo = 8'h8;
            166: spo = 8'h9;
            167: spo = 8'h9;
            168: spo = 8'h9;
            169: spo = 8'h9;
            170: spo = 8'h8;
            171: spo = 8'h6;
            172: spo = 8'h5;
            173: spo = 8'h4;
            174: spo = 8'h2;
            175: spo = 8'h2;
            176: spo = 8'h1;
            177: spo = 8'h2;
            178: spo = 8'h3;
            179: spo = 8'h4;
            180: spo = 8'h5;
            181: spo = 8'h6;
            182: spo = 8'h7;
            183: spo = 8'h8;
            184: spo = 8'h8;
            185: spo = 8'h7;
            186: spo = 8'h6;
            187: spo = 8'h5;
            188: spo = 8'h4;
            189: spo = 8'h3;
            190: spo = 8'h2;
            191: spo = 8'h1;
            192: spo = 8'h1;
            193: spo = 8'h2;
            194: spo = 8'h2;
            195: spo = 8'h3;
            196: spo = 8'h4;
            197: spo = 8'h5;
            198: spo = 8'h6;
            199: spo = 8'h6;
            200: spo = 8'h6;
            201: spo = 8'h6;
            202: spo = 8'h5;
            203: spo = 8'h4;
            204: spo = 8'h3;
            205: spo = 8'h2;
            206: spo = 8'h2;
            207: spo = 8'h1;
            208: spo = 8'h1;
            209: spo = 8'h1;
            210: spo = 8'h2;
            211: spo = 8'h2;
            212: spo = 8'h3;
            213: spo = 8'h4;
            214: spo = 8'h4;
            215: spo = 8'h4;
            216: spo = 8'h4;
            217: spo = 8'h4;
            218: spo = 8'h4;
            219: spo = 8'h3;
            220: spo = 8'h2;
            221: spo = 8'h2;
            222: spo = 8'h1;
            223: spo = 8'h1;
            224: spo = 8'h1;
            225: spo = 8'h1;
            226: spo = 8'h1;
            227: spo = 8'h2;
            228: spo = 8'h2;
            229: spo = 8'h2;
            230: spo = 8'h3;
            231: spo = 8'h3;
            232: spo = 8'h3;
            233: spo = 8'h3;
            234: spo = 8'h2;
            235: spo = 8'h2;
            236: spo = 8'h2;
            237: spo = 8'h1;
            238: spo = 8'h1;
            239: spo = 8'h1;
            240: spo = 8'h0;
            241: spo = 8'h1;
            242: spo = 8'h1;
            243: spo = 8'h1;
            244: spo = 8'h1;
            245: spo = 8'h2;
            246: spo = 8'h2;
            247: spo = 8'h2;
            248: spo = 8'h2;
            249: spo = 8'h2;
            250: spo = 8'h2;
            251: spo = 8'h1;
            252: spo = 8'h1;
            253: spo = 8'h1;
            254: spo = 8'h1;
            255: spo = 8'h0;
            default: spo = 8'h0;
		endcase
	end
endmodule