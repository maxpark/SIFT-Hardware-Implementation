.box 1 RISCV_P1_TOP_ipc_adder_8 17 9
.input 1 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7]
.output 1 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7]
.delay 1
900	800	700	600	500	400	300	200	800	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	300	400	300	200	-	-	-	-	-	
500	400	300	200	-	-	-	-	400	500	400	300	200	-	-	-	-	
600	500	400	300	200	-	-	-	500	600	500	400	300	200	-	-	-	
700	600	500	400	300	200	-	-	600	700	600	500	400	300	200	-	-	
800	700	600	500	400	300	200	-	700	800	700	600	500	400	300	200	-	
900	800	700	600	500	400	300	200	800	900	800	700	600	500	400	300	200	


.box 2 RISCV_P1_TOP_ipc_adder_32 65 33
.input 2 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CA[15] CA[16] CA[17] CA[18] CA[19] CA[20] CA[21] CA[22] CA[23] CA[24] CA[25] CA[26] CA[27] CA[28] CA[29] CA[30] CA[31] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14] DX[15] DX[16] DX[17] DX[18] DX[19] DX[20] DX[21] DX[22] DX[23] DX[24] DX[25] DX[26] DX[27] DX[28] DX[29] DX[30] DX[31]
.output 2 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14] SUM[15] SUM[16] SUM[17] SUM[18] SUM[19] SUM[20] SUM[21] SUM[22] SUM[23] SUM[24] SUM[25] SUM[26] SUM[27] SUM[28] SUM[29] SUM[30] SUM[31]
.delay 2
3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	3200	3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1400	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1500	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1600	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1700	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1800	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	1900	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	
2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	2000	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	
2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	2100	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	
2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	2200	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	
2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	2300	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	
2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	2400	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	
2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	2500	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	
2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	2600	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	
2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	2700	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	
2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	2800	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	
3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	2900	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	
3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	3000	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	
3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	3100	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	
3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	3200	3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 3 RISCV_P1_TOP_ipc_adder_16 33 17
.input 3 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CA[15] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14] DX[15]
.output 3 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14] SUM[15]
.delay 3
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1600	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1400	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1500	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1600	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 4 RISCV_P1_TOP_ipc_adder_10 21 11
.input 4 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9]
.output 4 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9]
.delay 4
1100	1000	900	800	700	600	500	400	300	200	1000	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	700	800	700	600	500	400	300	200	-	-	-	
900	800	700	600	500	400	300	200	-	-	800	900	800	700	600	500	400	300	200	-	-	
1000	900	800	700	600	500	400	300	200	-	900	1000	900	800	700	600	500	400	300	200	-	
1100	1000	900	800	700	600	500	400	300	200	1000	1100	1000	900	800	700	600	500	400	300	200	


.box 5 RISCV_P1_TOP_ipc_adder_11 23 12
.input 5 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10]
.output 5 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10]
.delay 5
1200	1100	1000	900	800	700	600	500	400	300	200	1100	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	
1200	1100	1000	900	800	700	600	500	400	300	200	1100	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 6 RISCV_P1_TOP_ipc_adder_14 29 15
.input 6 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13]
.output 6 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13]
.delay 6
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1400	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1400	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 7 RISCV_P1_TOP_ipc_adder_15 31 16
.input 7 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14]
.output 7 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14]
.delay 7
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1500	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1400	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1500	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 8 RISCV_P1_TOP_ipc_adder_18 37 19
.input 8 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CA[15] CA[16] CA[17] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14] DX[15] DX[16] DX[17]
.output 8 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14] SUM[15] SUM[16] SUM[17]
.delay 8
1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1800	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1400	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1500	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1600	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	
1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1700	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	
1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1800	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 9 RISCV_P1_TOP_ipc_adder_19 39 20
.input 9 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CA[15] CA[16] CA[17] CA[18] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14] DX[15] DX[16] DX[17] DX[18]
.output 9 CO SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14] SUM[15] SUM[16] SUM[17] SUM[18]
.delay 9
2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1900	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	200	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	300	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	400	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	500	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	600	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	700	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	800	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	900	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	1000	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	1100	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	1200	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	1300	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	1400	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1500	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1600	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	
1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1700	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	
1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1800	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	
2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1900	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


