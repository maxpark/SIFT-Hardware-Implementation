module HME_VEX_SOC_V1 (
    input               core_clk,
    input               core_reset,
    input               memory_clk,
	input               debounce_clk,
    output              memory_reset_out,
    output              uart0_txd,
    input               uart0_rxd,
    input      [31:0]   gpio_in,
    output     [31:0]   gpio_out_en,
    output     [31:0]   gpio_out, 
    output              spi0_clk,
    input               spi0_miso,
	output              spi0_mosi,
	output     [7:0]    spi0_scl, 
    inout               i2c0_sda,
    inout               i2c0_scl,
    output     [15:0]   apb_paddr_s0,
    output     [0:0]    apb_psel_s0,
    output              apb_penable_s0,
    input               apb_pready_s0,
    output              apb_pwrite_s0,
    output     [31:0]   apb_pwdata_s0,
    input      [31:0]   apb_prdata_s0,
    input               apb_perror_s0,	
    output     [15:0]   apb_paddr_s1,
    output     [0:0]    apb_psel_s1,
    output              apb_penable_s1,
    input               apb_pready_s1,
    output              apb_pwrite_s1,
    output     [31:0]   apb_pwdata_s1,
    input      [31:0]   apb_prdata_s1,
    input               apb_perror_s1,
    input               apb_dev_intr,
    output              sys_reset_out,
    input               jtag_tms,
    input               jtag_tdi,
    output              jtag_tdo,
    input               jtag_tck,
    output              ddr_port_arw_valid,
    input               ddr_port_arw_ready,
    output     [31:0]   ddr_port_arw_addr,
    output     [7:0]    ddr_port_arw_id,
    output     [3:0]    ddr_port_arw_region,
    output     [7:0]    ddr_port_arw_len,
    output     [2:0]    ddr_port_arw_size,
    output     [1:0]    ddr_port_arw_burst,
    output     [0:0]    ddr_port_arw_lock,
    output     [3:0]    ddr_port_arw_cache,
    output     [3:0]    ddr_port_arw_qos,
    output     [2:0]    ddr_port_arw_prot,
    output              ddr_port_arw_write,
    output              ddr_port_w_valid,
    input               ddr_port_w_ready,
    output     [127:0]  ddr_port_w_data,
    output     [15:0]   ddr_port_w_strb,
    output              ddr_port_w_last,
    input               ddr_port_b_valid,
    output              ddr_port_b_ready,
    input      [7:0]    ddr_port_b_id,
    input      [1:0]    ddr_port_b_resp,
    input               ddr_port_r_valid,
    output              ddr_port_r_ready,
    input      [127:0]  ddr_port_r_data,
    input      [7:0]    ddr_port_r_id,
    input      [1:0]    ddr_port_r_resp,
    input               ddr_port_r_last,
    output     [7:0]    ddr_port_w_id,
    input               ddr_mast0_aw_valid,
    output              ddr_mast0_aw_ready,
    input      [31:0]   ddr_mast0_aw_addr,
    input      [3:0]    ddr_mast0_aw_id,
    input      [3:0]    ddr_mast0_aw_region,
    input      [7:0]    ddr_mast0_aw_len,
    input      [2:0]    ddr_mast0_aw_size,
    input      [1:0]    ddr_mast0_aw_burst,
    input      [0:0]    ddr_mast0_aw_lock,
    input      [3:0]    ddr_mast0_aw_cache,
    input      [3:0]    ddr_mast0_aw_qos,
    input      [2:0]    ddr_mast0_aw_prot,
    input               ddr_mast0_w_valid,
    output              ddr_mast0_w_ready,
    input      [31:0]   ddr_mast0_w_data,
    input      [3:0]    ddr_mast0_w_strb,
    input               ddr_mast0_w_last,
    output              ddr_mast0_b_valid,
    input               ddr_mast0_b_ready,
    output     [3:0]    ddr_mast0_b_id,
    output     [1:0]    ddr_mast0_b_resp,
    input               ddr_mast0_ar_valid,
    output              ddr_mast0_ar_ready,
    input      [31:0]   ddr_mast0_ar_addr,
    input      [3:0]    ddr_mast0_ar_id,
    input      [3:0]    ddr_mast0_ar_region,
    input      [7:0]    ddr_mast0_ar_len,
    input      [2:0]    ddr_mast0_ar_size,
    input      [1:0]    ddr_mast0_ar_burst,
    input      [0:0]    ddr_mast0_ar_lock,
    input      [3:0]    ddr_mast0_ar_cache,
    input      [3:0]    ddr_mast0_ar_qos,
    input      [2:0]    ddr_mast0_ar_prot,
    output              ddr_mast0_r_valid,
    input               ddr_mast0_r_ready,
    output     [31:0]   ddr_mast0_r_data,
    output     [3:0]    ddr_mast0_r_id,
    output     [1:0]    ddr_mast0_r_resp,
    output              ddr_mast0_r_last,
    input               ddr_mast0_clk,
    output              ddr_mast0_reset,
    output              axi_s_awvalid,
    input               axi_s_awready,
    output     [31:0]   axi_s_awaddr,
    output     [7:0]    axi_s_awid,
    output     [3:0]    axi_s_awregion,
    output     [7:0]    axi_s_awlen,
    output     [2:0]    axi_s_awsize,
    output     [1:0]    axi_s_awburst,
    output     [0:0]    axi_s_awlock,
    output     [3:0]    axi_s_awcache,
    output     [3:0]    axi_s_awqos,
    output     [2:0]    axi_s_awprot,
    output              axi_s_wvalid,
    input               axi_s_wready,
    output     [31:0]   axi_s_wdata,
    output     [3:0]    axi_s_wstrb,
    output              axi_s_wlast,
    input               axi_s_bvalid,
    output              axi_s_bready,
    input      [7:0]    axi_s_bid,
    input      [1:0]    axi_s_bresp,
    output              axi_s_arvalid,
    input               axi_s_arready,
    output     [31:0]   axi_s_araddr,
    output     [7:0]    axi_s_arid,
    output     [3:0]    axi_s_arregion,
    output     [7:0]    axi_s_arlen,
    output     [2:0]    axi_s_arsize,
    output     [1:0]    axi_s_arburst,
    output     [0:0]    axi_s_arlock,
    output     [3:0]    axi_s_arcache,
    output     [3:0]    axi_s_arqos,
    output     [2:0]    axi_s_arprot,
    input               axi_s_rvalid,
    output              axi_s_rready,
    input      [31:0]   axi_s_rdata,
    input      [7:0]    axi_s_rid,
    input      [1:0]    axi_s_rresp,
    input               axi_s_rlast,
    input               axi_dev_intr
);
`pragma protect begin_protected
`pragma protect version=4
`pragma protect vendor="Hercules Microelectronics"
`pragma protect email="supports@hercules-micro.com"
`pragma protect data_method="AES128-CBC"
`pragma protect data_encode="Base64"
`pragma protect key_method="RSA"
`pragma protect key_encode="Base64"
`pragma protect data_line_size=96
`pragma protect key_block
UZud4f7B6/v6FxQKhmjyaTXeERXzfRip6ZtSNUmhYUG0Ald0RaoTpODL1JiArzr6R6R+9E0N3i80ZYIyD6X0MQAQsE4n3u82S73PXRVpYZgdax2PuWHX19NDCnfHaMwlHZhk6rVibz6pETkc1YTQtueXqZ+GM9n8FpDJcqc1fyQ=
`pragma protect data_block
rZY+XdSkH4lY6omSSWNTV/wsWsHHVj9HFditlIj96SJHbE8R0jHvFGkRAPbPyPGBSOcGTfEVDEsmsChfTGZ09EImvW9m8C0q9riVNVPk5buiyfutJRbFcmsdUT0jYq69
Qia9b2bwLSr2uJU1U+Tlu+3DoasjKp7F4ygMd5X9ipwdrE6KkQJYcNPPGXMfT6fIxECusEpiFSnG+v/qBVbVtJo9AVCc+bcfZYNRhmpMEfPoS9drRkk7n8ob8Tiw1zgv
rOQXrB+v79RvN9LzilLrKSlAaXXAP2T6ah7hoXNchzUBms7U/1rqrECI8pulTzrIq4AH5OudOyWNnCrJYzj5n6HD7gHgNvCFHg08idy36GbCeGlVO/DCgmv9+0YTEOIT
hMIpVq1eX7VMjnSHahnLCJDdT2rcUC5+gEQ/BhhH+/XNGqzrwixcSTbAr0elnZo58n6IGop6xjHO3cX05GH8xA0qN1s/lkaGJ7mGVPFgt49CJr1vZvAtKva4lTVT5OW7
MhvhoVZDLn9sFOCdyuyIcod0kaXgN0hJdI0qF4ITKnawrv3jvkttV1p4ZjzfLsbVPMWgHPM2upmTpyiyqCi8N97YN+iWSI0zfA+1UPUf1bLMPi04yDykY0/yz/RBIfNa
rZY+XdSkH4lY6omSSWNTV8s5nZymxHQyIIx3IqIdPAFY66gqgTFjv6CfP2dPNGWfAPz7zyDtY9nR+dtDYcf6iUImvW9m8C0q9riVNVPk5bsyG+GhVkMuf2wU4J3K7Ihy
W64Avqs5YPi2ZFOPEg79JquAB+TrnTsljZwqyWM4+Z9q7YBL5YrAylNP5/K6QVisR2xPEdIx7xRpEQD2z8jxgf9kcVp6zD5AMmeFX8QKZM0v2d4MiEeBQIhwDprEoW9H
kN1PatxQLn6ARD8GGEf79QJ+prAsJz4QdSNRq8crvNYFgnd7putLqzaUKlsbxcSst71fFIgTDTU9g1tTXr6k/d6J3SIBUl7FIzj0pH2Cva6Q3U9q3FAufoBEPwYYR/v1
An6msCwnPhB1I1Grxyu81vA8oG/pceRQxMUZCMLOS9wYqnvduVXPdRTHE+zwli3mguAq7H0tCd1HvLZdlpor5sG8nnWZcDRH+vdnptfcdcXKhutP56KtseqsBQIPMSVz
4o6UM47Mi6q7NI+YP+HQHU2kharRRGb26wS0y+Y2cGDCeGlVO/DCgmv9+0YTEOITqHd69sei06hDhJqIIln8uM4FdsQczP9JZb6SFGpc/WiQ3U9q3FAufoBEPwYYR/v1
uJg0Wx2RJWr5CTghvXzqpmd/+DKDaONwv4BB2Jg/3DeTKM1u+2Wg4xOxaWGRQL5Keus0wk8eb950U0F0gmaqZyfsXt9DfKq8UFD4F6nD5H+BIRQGKEmnt9CNoBbHPULy
eus0wk8eb950U0F0gmaqZ8+WYeFviGVKeqC2dk8krz3KiCbRJr2HgYyrX3ljAm2I74oAfe8PdZ0LQTtARvmiAsBCxI4pQu+Utgm/5t2LTMd0wYg2RvYn/PAGNKEI5xXG
Cy3A9C82rzhlol/lvapW8ZF0zGUPIeb7bWQasoaxp07Qv+fBbiZ7ZmTHPL8BJJgAvmQ/lT2dYCsEpsGArugKT/oiFHqHLUjtUhhvqeAmOo3Qv+fBbiZ7ZmTHPL8BJJgA
byeJOT7uu4H9ZaVnbdlqHrSi42CibOM+/jEPGNo3WyORKnzlGPAXWqgXZgRBSpt8BtdOL4TocPqFA/um7KGrRoEhFAYoSae30I2gFsc9QvKfZvX8CFkkHAn/NCRAIuEi
1+zFPsv/ySfgPsdtxX4vrsJ4aVU78MKCa/37RhMQ4hMxi9Os4c4s+ro/WecNNAfOIIzqwsZOs4cI+wabBS8q3D8FKm5rPSVoUcxXDk98C8ONn8yVzOJ+L2fQiC4XaSwo
rZY+XdSkH4lY6omSSWNTV12tjpoO2OV0mPf5nZ7Ym314KLBM7H/AxxyG/jk50+8Uafcf01YpHTUfhdSkhBxEmFGVszD9X9C7BdRzTSpglc7aL0PMVzjJWsEC7AJ7R1Lu
23iajBCwgP/c5j++AtTIa1JQqR+1W4klLyJKpPv1BrVriUw65Bu8J8OsNSP6bflqJIp7G/f7DpentpgqiX2Y7tm78p4ukCX0XZRhaDCO4fKLMtawqsVo5gs3KrDV0oap
mWw1ojcQcdc8Ty24t41JnsJ4aVU78MKCa/37RhMQ4hOBf1mIweWhlVpijFiWuvTjoF2lhZBrJBUmtVJgOTOm8ZDdT2rcUC5+gEQ/BhhH+/VA2OOGMwPfY31dQsL1LAb4
tHSHQXWCzus3ROdc345RXnc2EUmKaxFqwQAYeiKQNUehO8/whGWZxYm8jo2M/dFc9gqliS9njW5DP7ndTCUT+pgVy4OxUdW8OdbLX0G3Sj2mw6ef9G/a9tONSX+UVixf
EZcr6lMAtC68qySmbf2y6lGfKvss99kkAFlBAcwKnwZgKPmihm1usyNCx+mcwvln+l0Q1885OqRM8ejd6UbkkQrjUhoIMMVclD6PUVEARytaL6r9Dmn23DcuArBNiH6y
+l0Q1885OqRM8ejd6UbkkarMxB7T8oZSKJ3kwyGrex3HidyUqTucTGyXOUsShleEHgPg1mwgPBDqhRwRuQJycSVqm4W4iUIAf6opdGDLctTld83jZdWZezTgECU4HnQB
sjdB4BBS8+QYihSzjty8XZF0zGUPIeb7bWQasoaxp06wg2pOoE8zu82q87VU0rayv0qL23AYWi5UAsJ0luGLHvhhO0TE28YpxF6+yBua85VSaM3YW+iOYEhTngayst1r
14+BkIz7OUtZhU7l2s+Kkz+lH6IAuvCLxnvcVy47fbd0wYg2RvYn/PAGNKEI5xXGxUZ3Swg2+FQv+HRHg3lmYBvpIh0XGlq3WRwyhtYRMRmtlj5d1KQfiVjqiZJJY1NX
VbgSpfPCUUD/OTMLf1R6tKEX/inInUbnztgmAyvsmUPbeJqMELCA/9zmP74C1MhrnVM0pAtNJorVwBRAL2Qvkjrdm7vKdpOmhArfBDpzSKmQieSRPmDxdNsR9S2zblAq
sY0fvbSNx0+MJqfNjmpwSdu6+LDvqdi+9PkQxQs4MvI63Zu7ynaTpoQK3wQ6c0ipA/1sSabum0a5+IQ7CMWTSvd8WKW1IN/vgTHI9m5zwE4p8KMBcX/e4EporiZb4/0/
OPsJ6yHEbueMn+7BSrjxMcakdCWPm8GRN5J2SM4b+JKf+GkfYiIalMywY3yWE+3vmHe529OTjppeeWYxjDul6ZFCiwh1IuqgR0pyWBMwfnIxYmf9TfvieZq4i1+4laBe
gg3yWeL8eajASjlxWTSoVofi37CEzPd2G6nTl+T4wxr+WNCKwabbQzJjx+iJHz5ojnv1eBojtsvOm38g6CRlD/bRkA6qx/FSm9WXbqPi3+bYM64+dvN2Pr4PzQ4z32/U
S22E4gg7fIlH6gNoFoJ0Mj4RWNyWGTkYxU2oagczuoISA7E9a3GbtWs+QQ36MbkXWu8oEzO1OkvbgY6SphNl6nk6Vp5DPXvakUvltpXQWm1/0KTxvCSFaxENyjQL8PhC
GKp73blVz3UUxxPs8JYt5pSJ6gOXAwDN3byP8PoQ1linAZie5JdVbbTv/pElS/YQkN1PatxQLn6ARD8GGEf79Xb5kkF2aAcAO9dv9SXXJUl/Bhr1p3ObmqB0MFqgvHyW
vbWNJY6eTH4cqDRKSZ2uQD1SS+WnWY022WBiHK1CLHpa7ygTM7U6S9uBjpKmE2XqaAoclGunj7FiEnNNNrZqj97YN+iWSI0zfA+1UPUf1bKGJ9Ma14fZ705U9Q2F/w8F
skgmMbaKurzT40ERGlWNLjFiZ/1N++J5mriLX7iVoF6Jha1wUIpMRUWKcuOz7vERwqVUWUUhjh9zeno38Os8UoCmNxzirTYd7fXcs4sXVISE3gtIYGDNgDcBqq8eNgMj
7L0y/1+Dc5NnTJtwm8+ATcKlVFlFIY4fc3p6N/DrPFLH7cWWtjqjHC2Y0vTybTd7uY5z/UiHUqwsHvmOrlepRNphABHXVkl+LUfoFzZj0kuh+RsMv0BamRMVKntu1hXl
yMktjPWKdmH0j7N80rEt/pDdT2rcUC5+gEQ/BhhH+/V2+ZJBdmgHADvXb/Ul1yVJCnNnEh3FzdTOATiHzbDWEtdIIG4OVopyISytWsbuR3YYqnvduVXPdRTHE+zwli3m
Ei4olFzwV9zmPES+X4ONMTGJmAjvDvCCPzVsI/eJt7C5jnP9SIdSrCwe+Y6uV6lE2mEAEddWSX4tR+gXNmPSS3BkeGBMQMtr94W7uZn8JsSApjcc4q02He313LOLF1SE
hN4LSGBgzYA3AaqvHjYDI+y9Mv9fg3OTZ0ybcJvPgE2H4t+whMz3dhup05fk+MMaZOPBketMLMQJFkuna2gtQfoiFHqHLUjtUhhvqeAmOo0ijse/2fluE1CGerRdUSsg
HvwXsbFdJGAcVA9TXeoOKCACg1ghTsA3A4l07RS3dJUCUeoWObcQ13BCzHrsHY2v74HCLaUerkqzF3L7n3b27FrvKBMztTpL24GOkqYTZep5OlaeQz172pFL5baV0Fpt
UZ8q+yz32SQAWUEBzAqfBlu0YppEZjnLxDzROYLlq71a7ygTM7U6S9uBjpKmE2XqeTpWnkM9e9qRS+W2ldBabbMZz5ULbCOlbZsFhAwb+PlCpkhNV+qPCe4K76e1jad0
Wu8oEzO1OkvbgY6SphNl6nk6Vp5DPXvakUvltpXQWm2kw72h0yEkAQK7hrMsWNsxdMGINkb2J/zwBjShCOcVxh/HklvYg1eOzX5kYPaydni7oqcFMPW1kp3UhB5HeLTC
KkHTYLZ3eFVgR6Fcq8b8rDeWEXXDgUAgj9Brh/+atheEM4JIbbqrqQcYanvjF2CegAdXtwqDtrkMcTULh34OFBKEqu5eY4moQkLgYLOWYjI5kiYzkhCpaaVJNvC8ms5K
G30DxeGu1xUPnxN/RXzT/K2WPl3UpB+JWOqJkkljU1ekW90qF7QeuvFSNZKPUlveBONagr2PcZ9zXBKBZWw6OZDqAv8LbHKLlrhNYS91Ol0U+u2gQq5qg4cvhJh99JOn
HNfuQvYsDCb1r0BdkJ0NGsc40kxf+lZn34bO1gpWUTs8NN25+d7Em112fBjs8rzJ/63B5bY+V3O5Dz9xYiPHkoCtrRvQiix+8+hfsyuorTpmLNVzb+wDcWnY41obtPJp
g3+pG+FbCO8oTTvnmsqw6xT67aBCrmqDhy+EmH30k6cc1+5C9iwMJvWvQF2QnQ0aq6eKiSKExQyid+sIBxb1y33NKbyn1fO4kh+TP5E9N7mALFP3rF4vLbSjTQHuSXxR
rZAVMJhttom2tDl6Mt0nTbuZSQuv2LYCQq0qfBr/yTlHbE8R0jHvFGkRAPbPyPGB0Z9Vd/k3UPnD1WwwWCRXPpQW1p+rm+iQFPAWFiwbNWvtyUsOJD3CS85a7SzIsCE7
lNhXxYsj+33nrPEXJNnKOBzX7kL2LAwm9a9AXZCdDRoaqt0T08p//ag3WizGQaDsi5IpdFCcD+FVTbzsNb9+2QDHcaR9oXg0UaSnAcEGw2HosGB6pZQdm+1gU+V2y25p
SpQjZhGRlVE/MEN0103Z71EN0XFVS7qPH/APwydBTrEVTIXp1esBpr7sFht7fqFXCmG8PVkc/R3SGqZJPSgjDppHonl7MnRuBJK4DkzTLxGLkil0UJwP4VVNvOw1v37Z
AMdxpH2heDRRpKcBwQbDYeiwYHqllB2b7WBT5XbLbmnB1gGZ2R2YveulqOgjblIgwnhpVTvwwoJr/ftGExDiE7elb0EVn49vmGinvJqr9pfWXINnDRtRiKbGz46nq5RW
afcf01YpHTUfhdSkhBxEmCUCDevj9DjJ7PA6KtyYmSD9LnbcR/HHCVRmbWznPpBePFVS5qefGUCjDRjqZ5IvdH9FVK2W5QmhsFNwzvOAkmKj668iJj8ZicsD+lHn5taU
sqy3gzfS/Ab7LSu1771xb73N6eugI9QosBXhV4l4rH4U+u2gQq5qg4cvhJh99JOnGppd/bk1b+rV99JUv7QLv3wBsaKbAXC+3OGiD5pfLhqxjR+9tI3HT4wmp82OanBJ
464o4j6QWBRQLQ+usy+Meor1y528GyE0wZFn88jZ4bNk48GR60wsxAkWS6draC1B+iIUeoctSO1SGG+p4CY6jTBl84EvpHCRbjrqj8nYeYiK9cudvBshNMGRZ/PI2eGz
n/klliVLMhZ5RiAytKoqtMMBfzJZ+Jt6QrfNPqnQBGLJ9UQPF/dwtZ0w3z1dXKLwAoXMC4K/9xP/SWOt6wzZINv5AiHFH1vvyi0kUwhdOmOwz6ws4LfIaOjE8aAGj72J
wH1AWcP5taswW+0xmqVgvs75ZK4RrN0XbAjOBuhrJRRlYNgUgDVcEjiOk+iVgCyiT4o+ycFjNLai+e5fFZWDz7elb0EVn49vmGinvJqr9pcbfihAz7uVEbgyCGk4GuBc
wdYBmdkdmL3rpajoI25SIMJ4aVU78MKCa/37RhMQ4hO3pW9BFZ+Pb5hop7yaq/aXhunPfztBF00NP3VNuuzCHw8kxWRPpKAatSVRsRjAsz8NvUIyoebTorkGAdMF5EJD
u0A7EV1bdj0SoV9IymjICF/PzRQgublauU/DapG9Ts8PJMVkT6SgGrUlUbEYwLM/Db1CMqHm06K5BgHTBeRCQ7tAOxFdW3Y9EqFfSMpoyAj0pvrJI05RhDQJ9zN1zKja
afcf01YpHTUfhdSkhBxEmA29QjKh5tOiuQYB0wXkQkO7QDsRXVt2PRKhX0jKaMgI5Kz9ntvELDvWF3pMyKCz3zFiZ/1N++J5mriLX7iVoF7SBoIDIgS70Hh3ir23GaAv
HtJLa4LCBk/QpJrL5CdRIY3WUseYTOJjnm586pqEQkwfV4GzoqgfXIVSWNJUiXTW41FnfCeZkFJmaJwalVa5hAqJrloSNP0zFCLM92m3MQDpihAanr3fh1KE+ukRthhF
10+KIXsFYTOG6b0aut2at08VkE5SNQvAY1Mih8waGeKD9KhGbwWqAGk+9B3WFPLOAuocZcRiEJ9sgcbvLV3atqty7OMtbsWm+GIZn/WPh9061clngAlWUiSuYbTFMv8e
R2xPEdIx7xRpEQD2z8jxgcxWQSoulk6kcHsQHzLCmXA0sTxSc3Fb+JQMAdAnjo/Jvh198dSkCdiNenzlHMVWs5MozW77ZaDjE7FpYZFAvkrMVkEqLpZOpHB7EB8ywplw
NLE8UnNxW/iUDAHQJ46Pyd9ahynKKek20ZVTZFeEA9/oXK2y2IwAlLo4rGziyzxIXoCllUOkzU3SH8hn7OXoEW0xohjSzRs8thLEX+w+oH9XehkbOBtSN0BkfU3yye5n
kH+R5iaAROlsVfKBgS07agqJrloSNP0zFCLM92m3MQCHz51KHGIS3SUHm6DHEstpZtonhaiqZp9i24j6pCrwnLr/d6zTt+cL7zyOVXqI7NDkitwaGdT73c2EeXEwimmy
CzA1giAT9fiKUkIvtLOxqhWhRETpFpmMz2OGYFUphWQbrxcGe7he+qeufjGLZjeI5IrcGhnU+93NhHlxMIppsgswNYIgE/X4ilJCL7SzsarBZGZkZAZ96aFHtwj9i+eh
5MTHwCPNcns/aMRXjDbE3p1flbsnOLtaHTyQKADNnOq0X6/E/aDXWfbBZX4t1noL4UHyxb4jyKK13WkSWdYgBeTEx8AjzXJ7P2jEV4w2xN6dX5W7Jzi7Wh08kCgAzZzq
WVjmuB5r0rI62RBLMRyRXmj8ewgqg9dlJQPyPPXvxdZcamTE59vtVchwulaqZIfByHfX90Etu+C/RxWSmaPQ8vnmzcXYi9xLwvLlzYY8oE0PJn96Fxr7rt7ZrLcbKE/R
KOU8C4/a+ylMTlwuCQYe+zpFaV9ZjyW0vKCFXl3gH2/xONENfwAq8j+cXrJiQZg5KkHTYLZ3eFVgR6Fcq8b8rJ80Bi6sypPV30l0Oewc6hse0ktrgsIGT9CkmsvkJ1Eh
w+/7ZNvs4gSGSkEpwQNOfkdsTxHSMe8UaREA9s/I8YHMVkEqLpZOpHB7EB8ywplwNLE8UnNxW/iUDAHQJ46PySUc7mq/UkHm79iScU28h9je2DfolkiNM3wPtVD1H9Wy
3cNOtmIzWwWRh9hdGn3AGCAHxV4w42/CGkuvd/kkXcZYoW/Fszry4r0JGDFQPDXG3A/PxgQYWgYJCytdn1VqUT0wjltC+rQNEVP1Kn/fNi5AEgRC0FyJT36UXLOSPS0s
5WETENxKuPyiLnikTfu9e+TEx8AjzXJ7P2jEV4w2xN7SBoqsTXZBfKS4CqWNm/17F9QXUdJt4JdO9U110Sgc4L21jSWOnkx+HKg0SkmdrkDR5ShRIl94UvBsC1M5FJnJ
tpzsxfRgVAH0LvQCU/Sx14PM7aVoqS74jNuQs2qA23W9j4b+2WyrQpbTopmuMgK6siOeRKBCBKJAzYw1Ewm/eTRi6/Q7+mjbCiqWtUGmNqxGTwhAhTqJySTqaHKh4Fuu
ad5aNGtSdIRM8ti1U/N7qFA6uSfJWcRYAvcWI279ogCHWZVFN1C4ZdsqpdxEhvEcdeNnc0aOhiJ4MScrISs9raYrXr2XWga/PP8eqyhYn1jkxMfAI81yez9oxFeMNsTe
0gaKrE12QXykuAqljZv9e8+nuuQS4tsf30Z1z9sarxYK41IaCDDFXJQ+j1FRAEcrVUxXCTVmMrFaR7Ru5Hr6hrac7MX0YFQB9C70AlP0sdf1Njtv6wj3oZ77RtKPrE8V
QE095xHecGbrNUtbeCSupUgYkj1yTntkFNGBfPjz/LV9RShOX4pAd5/GmofNusGvL/TrlKgUdFkC0Kwq+Cinc7scyheMGBf297+1s5w5SCOveyi0N13qZ4pHIXwmOETs
CaqiCCbbB/U4/0qxioQZGw2bvtGZ43uxx517P/doAvOAFRcKFBbiOT1X/jSJQtiN/6rmdjtYG/ZLKsscErsBSH7TlYSxBg1zyS/566rxLvnbeJqMELCA/9zmP74C1Mhr
67CtcLqZhKaAsp8/23T0oNZA3k0EnrdhFInzGNbJ/NwdiIojrXJTEu1goQstByaYvY+G/tlsq0KW06KZrjICunREBWtlKsYoCp6biz44K5w0Yuv0O/po2woqlrVBpjas
0G86My8ur2VQJ61XLMVkFuzzOnG81fWaUX2+9m5kxvf/FfnKlwuDhGkgzE9MBMdsZ3JCNYv2zsw6O4Y3Fh11p420BXjy3fAxMTfcc0c+NzgKDLQ0qQCNovUuexI/JyB5
4vxlw9YuKkvFwCnfglX19g5pQuUrhjkblzQeOns6JP4Pq4BOhJj1G/UDo9KKqvWk6FytstiMAJS6OKxs4ss8SOL8ZcPWLipLxcAp34JV9fYOaULlK4Y5G5c0Hjp7OiT+
BUb9eRfA1fUpGVYL8hfg6huvFwZ7uF76p65+MYtmN4g9MI5bQvq0DRFT9Sp/3zYuaY3SecHz2Z+yApnqIuEE+LJ3FPmhMbQUy8qeUDvCBUQxLFNhjd3n4e2W74alQGlS
/6rmdjtYG/ZLKsscErsBSEjWaHUU0KHyG0OFScn+mBlwO/BIrUnSQIyc09k3kZ03GTZhDcdAs/G6pfDxOz6WYZGlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKU
p6lR876yb+Qf7IBKwJwXeN2PnuGEzA48mYnK/iSbVh+HWZVFN1C4ZdsqpdxEhvEcjjVPZKIzjxKIDHAzwjcYBs2fupGwogWYqFQ9xxh5mm0o3uTf/NrlvMExTlVbTVNW
1kDeTQSet2EUifMY1sn83BZl1CGUpljS1UCH4K1fvIV/FwudDKXKnFmdEuYD3eGw/xX5ypcLg4RpIMxPTATHbGdyQjWL9s7MOjuGNxYddaePT85aSz46SLmj3xEKOrkV
rZY+XdSkH4lY6omSSWNTVwcz/AzImCCIvXvC41biajt1wLoUYjnAAEjwaCBgCZ6KzrkTQcKRUsbNbsSmexFwDEdsTxHSMe8UaREA9s/I8YHhzF75bxPWLnSIW6pOQxjQ
/1o8T2wfswjjZ88jh3VreR4H5PPAirs98ntcRbnyoHXjUWd8J5mQUmZonBqVVrmEq6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCHYfWOwu6JzilSG7DO4xaua
rxuXAPkhn4JZkRIi2C4K2JGlCOgXQweHAWpAKrw01tKwu9Kefezrr3TCcx3LMvedbnpoD2U1vqLsusnlUlwyy8oo2YfC5sH4iom1/1pAsmQ0Yuv0O/po2woqlrVBpjas
Oxsr/g3xgfx3jHvI4FrMSa2WPl3UpB+JWOqJkkljU1cHM/wMyJggiL17wuNW4mo7dcC6FGI5wABI8GggYAmeiiUc7mq/UkHm79iScU28h9je2DfolkiNM3wPtVD1H9Wy
r3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWfd83QsY7rSOy9S3cRsp9bE5MTHwCPNcns/aMRXjDbE3ou06eoRpvugoIqqlwLGYyn+k4AGmo1uZj2nWmBPbeMS
kN1PatxQLn6ARD8GGEf79fGIOR0z5ySwA+0bbOYvzYwxCHLrNnOQuZ3elaRhDK6n6+2BhyKwcO/WVVzDH3PYz8vvygXEb8unvqp/5eSvJQo2QxAEmEQ/TWxIGBuiZgrc
02yHNLjiqK7MNZflawE2V14zAoiHJVyWehBeVmBbqgbILWZQpoWgA32jr9HoBvFiyYXvFw1XoC2dSWCfoLIohx6tKuqEDos1vDoKMegWEpK2krJ9F/Tb/y0eoCrQ1m46
zUBH0P+b2ClmLFB+Gv9Csxy3g5OvxgmIWcSZjgnJreyQ3U9q3FAufoBEPwYYR/v18Yg5HTPnJLAD7Rts5i/NjJWOxeMm1rt4+c2ie5z3UvztyUsOJD3CS85a7SzIsCE7
wMMBAw0duLRDbA9vyI+EOTZDEASYRD9NbEgYG6JmCtyKJoTypdm7HSRqIc3qIi9Meg1ie9QNA0DUgSpBNOJ3zYu06eoRpvugoIqqlwLGYykmKRUT6bP2+AZJBzI9ZtFl
RMe0g7shdEuSAHNcBohXCc8oxwxhq9Ib5mKIG72IP9ulx5dViA0ouFLHDyJzCFRHrZY+XdSkH4lY6omSSWNTV0APjcsG5V+CsAumu/zdHmmjZGr+ga4/tRzeOFIPbGpB
qg7w03osV3q3/l2i+eboiMoo2YfC5sH4iom1/1pAsmRZOGFKjEONg3Js24m1eZiQ6zzsXpRNIxI6RaHrh0RcVdwPz8YEGFoGCQsrXZ9ValHILWZQpoWgA32jr9HoBvFi
Mkb7LYmLkkF3IOIBPMXsBq2WPl3UpB+JWOqJkkljU1dAD43LBuVfgrALprv83R5pYzrwpKjBQzz+BTh6iN1q+OP9uRzUEnHTeJuWizEiQUy5evGTaBq5M5mI2DxoC69r
caxCVjjDXntsopWrO2r2loxhBAIJmH9WJriaFqIvUzgoVHIKMbS+apsVZ6zCe/umRH/coTWKgENRZ0XCeml1EgfiU9p3WAaTsw/NaDHYc+tFYDecDkBvgZn+lEGu6OLC
3A/PxgQYWgYJCytdn1VqUcgtZlCmhaADfaOv0egG8WIZkGud0iRqu1bEcmqjetIF+KJVM0+aJm3SNUm7Jk03knjyxkGc/O/Cv7EBu412URmPfjSmrRhoK1/2nYH452YR
TxWQTlI1C8BjUyKHzBoZ4p2ZcrG0X+YmU1i5UdRGSFxZOGFKjEONg3Js24m1eZiQoeoYVEbkn4qi7/A2afXv4lA6uSfJWcRYAvcWI279ogA2QxAEmEQ/TWxIGBuiZgrc
gUovm+kYP8FZ8VoLRlBA6OTEx8AjzXJ7P2jEV4w2xN6LtOnqEab7oKCKqpcCxmMpsyXzL9eTGKca4UjQK4TEz8J4aVU78MKCa/37RhMQ4hM7yEf8Obx9sNllv8SVXJcL
vh198dSkCdiNenzlHMVWs5MozW77ZaDjE7FpYZFAvkrI9VqEMfWQG5zLG3renFgmW4aBGLSmyOVe85TZMYULilB/IRX200XvR4OPJtv+V8HI9VqEMfWQG5zLG3renFgm
LziblCRO93WJvIWH5+NN0Sc9TI8VVfxwqk77JJv5rcif57V5hGbPEjYgFY+1Auvm4hwCXIpgaUlbyZF9vvMd5lB/IRX200XvR4OPJtv+V8HI9VqEMfWQG5zLG3renFgm
coIDEA8qzPjg/wWbmFAS0x0OcNXhW9CWE6yq21HjWOY7yEf8Obx9sNllv8SVXJcLT667CVosQrbX+o7yPgpcDit4yzJRwMwbtPp+vPYF5BE7yEf8Obx9sNllv8SVXJcL
GBJxS5OJXvnZLZfKQssFXQ09ijq7E/YI8fcKPbpp0T/I9VqEMfWQG5zLG3renFgmJpFCy2lQbaN6vOqKcBlKkkLZJnxFLR+05+2wLmZ9l/vI9VqEMfWQG5zLG3renFgm
D0d5asSp0xqAZAeby1C1mmgjPa9L81g3aFJI8x56i+lAD43LBuVfgrALprv83R5p1KEJR9udbsPwZxDBD4GkgYEhFAYoSae30I2gFsc9QvLI9VqEMfWQG5zLG3renFgm
dNhUbvAYGLXxcutQMYS0P0dsTxHSMe8UaREA9s/I8YHI9VqEMfWQG5zLG3renFgmX1OlTvogl1uY5vvAfJBpr62WPl3UpB+JWOqJkkljU1dAD43LBuVfgrALprv83R5p
eiPZA7RRVI2iVqJyyZDOt98ctBV9iAOJmsnxuiIIJOZ40bc5fdGZ46VUz5N6wM/M9AVoU90rl9yHODlzYes4do9msKNMg75D69bo/5X2Ymqf57V5hGbPEjYgFY+1Auvm
tXXa5rnpwb/5HtSv+1oeYtwPz8YEGFoGCQsrXZ9ValFWNhi82WE/OvQ+gdQ7O2WUqaHdpDg5AfZRxSmh5fLsE4AVFwoUFuI5PVf+NIlC2I0sgVUgv/jYNp75ydmyHs99
tueDTG02eV391IQuObuPqZoGCa5kSQBKDk7N9B5yBebNtf/xkJR6UbxgwL2d/P8vvbWNJY6eTH4cqDRKSZ2uQNHlKFEiX3hS8GwLUzkUmcnvDGEAMYbloer5zJIZOvDD
mb8uiz9AxSX9ZtnfctfhteTEx8AjzXJ7P2jEV4w2xN7nIgz052WWswq9py7tYm8L8xXIL3kuNLnW4kvgxoGJ+7bng0xtNnld/dSELjm7j6maBgmuZEkASg5OzfQecgXm
T79jZcbf97PBlsoX4ec8sbyuxsjZgVDxPkAQzjpa6Kvr7YGHIrBw79ZVXMMfc9jPy+/KBcRvy6e+qn/l5K8lCmRcNwQ7ub5FuxILF2M1GMpmeZ0qCHzysK0SEVcLu+OL
DyTFZE+koBq1JVGxGMCzP8j+T5P8di6XieeA1YJl3frWjw+XAyK0VB0/bjMAmj0/VwkDJJ1sNFzsWZUm2mHIBAssUtpMXFjvdawCkkQSK4WPFW8f2WkNPKvmrCzQ8Taq
rizvr5OTPRaSaxKTOXKv8XyaGP+WdLegRtgA7h4GKSbmjYZGTPpx5fHkDH12aeTGU6bgO2hzpVM70iDAxRsbWz2UHhRP5OuAUuUz9JhC5sCh6hhURuSfiqLv8DZp9e/i
UDq5J8lZxFgC9xYjbv2iAGRcNwQ7ub5FuxILF2M1GMpDK4v/EpyPg+QzAIJ22PNNKkHTYLZ3eFVgR6Fcq8b8rA5ZwkuEkfiR8Ko9M3TERx1kQqy2K9YjZeCH1DEP2Kr+
gbuM4RHDh6Hq8g78wGEfPsJ4aVU78MKCa/37RhMQ4hMqNJI2EaH15panZ1qif+cJokiZvM70sM1kay/8QwD8u0pw6PAK/4tDiADewEe++KC6/3es07fnC+88jlV6iOzQ
RK6q0VoLiyzL4hM5mmYYxwnyKaneo3NdPxy6khV1/A8uovWMp1YmjJm2+98hLmZXuxzKF4wYF/b3v7WznDlII1Uh59ERS610z74PKFcPQirbhz7dQNpnag0SBmEdCDMe
HLeDk6/GCYhZxJmOCcmt7JDdT2rcUC5+gEQ/BhhH+/UEAryO2LIZOMoPRLzF2cA7KUQ4MOY8TOL4inlOOB2rQy4mPIfaZvE0zv8v1vTXUUCTKM1u+2Wg4xOxaWGRQL5K
SzWLLq88EuSCMnNbkzjOcX/hTbmkJA+DnpMVLDyIrXTmWxiTecsbiQca6IkQNSYt5o2GRkz6ceXx5Ax9dmnkxlOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4
w8pC2SqXiQ98WH/Q6n+MNewxYcfm5JQJ1VLe5bXzen0InAvfIjahchYT+82i/kG3OafClgp9xdeAiGEGzVGxiQD3KFCG7n2bV3zvfnWuw3ZBtXl17RcarRSYB7WlRBqj
ZFw3BDu5vkW7EgsXYzUYykzoN8Q2yYOgYPmjhaNy7s1/FwudDKXKnFmdEuYD3eGwsJBKNsb+RWp6tXGzrerfOWRCrLYr1iNl4IfUMQ/Yqv7PxDIyz+/dStSXxSVMGq4D
KFRyCjG0vmqbFWeswnv7pks1iy6vPBLkgjJzW5M4znF/4U25pCQPg56TFSw8iK10AV8hZvJ7UQYq50u36hzTPdJMZ45uzt8r0f/MToicFDlVIefREUutdM++DyhXD0Iq
3WH2CkwQjc8NjMfDzPFy6zzHe/YKIvDw+s8jrBszLWRsQlaQqXt+jNMreIPOEvi05yIM9OdllrMKvacu7WJvCwaG2BEPjYdOhFjTn0sB4mOrRU10XbAqFT2AH2j1tdBx
/ozHgkCqtaWGn4lSW4utgE+/Y2XG3/ezwZbKF+HnPLHkcXvBYihGAhgX7o2pMAFY+NuCJSqWsDli2Ssdw53wSGENuthXUW3WYQBD1AmUfHHgCA0O/fOXRBXvmcvYIB0R
pJm7IksAe4//Z1QoqrXw0JDdT2rcUC5+gEQ/BhhH+/UEAryO2LIZOMoPRLzF2cA7KUQ4MOY8TOL4inlOOB2rQ5gLM5whebiSqQ6KOHJs1E2TKM1u+2Wg4xOxaWGRQL5K
SzWLLq88EuSCMnNbkzjOcX/hTbmkJA+DnpMVLDyIrXSB3Fn6CSwc5UTqtQnvH+Hs5o2GRkz6ceXx5Ax9dmnkxlOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4
FMmQfEzPZEA34WSlrOMS7ewxYcfm5JQJ1VLe5bXzen0InAvfIjahchYT+82i/kG3iWBoDE8SXqHwT+E2TNJQLgD3KFCG7n2bV3zvfnWuw3ZBtXl17RcarRSYB7WlRBqj
ZFw3BDu5vkW7EgsXYzUYys+6OXEoqsLMu05Tkhok3vp/FwudDKXKnFmdEuYD3eGwsJBKNsb+RWp6tXGzrerfOWRCrLYr1iNl4IfUMQ/Yqv7x66PKvdRONz7kWa+US2Ac
KFRyCjG0vmqbFWeswnv7pks1iy6vPBLkgjJzW5M4znF/4U25pCQPg56TFSw8iK10aNupY3mzWblgmTS3JY75fdJMZ45uzt8r0f/MToicFDlVIefREUutdM++DyhXD0Iq
3WH2CkwQjc8NjMfDzPFy68Ym9pLWsEndRICWMK09ydRsQlaQqXt+jNMreIPOEvi05yIM9OdllrMKvacu7WJvC7w0GyVjq6iKYKfCB1NVisyrRU10XbAqFT2AH2j1tdBx
/ozHgkCqtaWGn4lSW4utgE+/Y2XG3/ezwZbKF+HnPLEAiqzfpuKYjNeBHpHzyvyy+NuCJSqWsDli2Ssdw53wSGENuthXUW3WYQBD1AmUfHHgCA0O/fOXRBXvmcvYIB0R
4Bea4M8GdLu4CCxKjod5i5DdT2rcUC5+gEQ/BhhH+/UEAryO2LIZOMoPRLzF2cA7KUQ4MOY8TOL4inlOOB2rQ3Vfu9ooXyVvntx0jaacivxW47D3lJA7/VDt8o9h9Auc
KjSSNhGh9eaWp2daon/nCaJImbzO9LDNZGsv/EMA/LvNJH+33d430cyIPrZOeXiCbEJWkKl7fozTK3iDzhL4tOciDPTnZZazCr2nLu1ibwvAnd2/OCubAlyrrCMXLGKq
67yBrpvrBP/q4kT/GpxqJcvvygXEb8unvqp/5eSvJQpkXDcEO7m+RbsSCxdjNRjKId20p1wMJ2gcq2dHcZluQypB02C2d3hVYEehXKvG/KwOWcJLhJH4kfCqPTN0xEcd
ZEKstivWI2Xgh9QxD9iq/kdE9efs0w6ga7Q2I/WJEOFHbE8R0jHvFGkRAPbPyPGBSzWLLq88EuSCMnNbkzjOcX/hTbmkJA+DnpMVLDyIrXSn/h1kNg1QFT46LQi8IBUf
yogm0Sa9h4GMq195YwJtiFOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLnT1QBVfdejt0d5UNJrNOblJDdT2rcUC5+gEQ/BhhH+/UEAryO2LIZOMoPRLzF2cA7
4NhFrwxGmyqHO+jR+TAV7Uz+/wVfV6Ukh1FUESF9lw3r7YGHIrBw79ZVXMMfc9jPy+/KBcRvy6e+qn/l5K8lCsDlicVnrgUWDK9VOIDcHDfvo0+10cUMbokuNWvWK1k4
n8B6Q5pOCez9vZLsayarneTEx8AjzXJ7P2jEV4w2xN7nIgz052WWswq9py7tYm8LlND94lvC14gXu5leKvPbMlyRAGy8PlAe92xJGRk/rQVW47D3lJA7/VDt8o9h9Auc
KjSSNhGh9eaWp2daon/nCQAjhmhAEFEe3H6UY3ibQy1l1nd9RnjgA8ls+Hk1EpjIsM+sLOC3yGjoxPGgBo+9iSr80b85AWN1ecJ1V7ghNmzg2EWvDEabKoc76NH5MBXt
2lV50Z8ZbO7R/XZAtMAgLOzzOnG81fWaUX2+9m5kxvewkEo2xv5Fanq1cbOt6t85/mXNNhQuNixZTrQ+ERII5Xfr0+zmQzh2JNUBLWruLao+7p7JGPm/+PG7fTw+hCvA
67CtcLqZhKaAsp8/23T0oNvqcSol8XG6fW5VWX77FzCfeyJXtRfpJuGzHxoBJqr2xuKs47xAlIb+nFZyvjXR6poGCa5kSQBKDk7N9B5yBeYEz7OH7NQB8S0bGD5jOdV7
qfefUfdWnFSGoL7piGzzIwqlIb3DfkHwCtidqYWxvDjmjYZGTPpx5fHkDH12aeTGU6bgO2hzpVM70iDAxRsbWxyLJM9m1+hZpHDVGPttMueInijiFB0YkuN03Rua0qMK
Hq0q6oQOizW8Ogox6BYSkraSsn0X9Nv/LR6gKtDWbjrb6nEqJfFxun1uVVl++xcwn3siV7UX6Sbhsx8aASaq9svCUc90x1uyyIqzT3Pxc1atlj5d1KQfiVjqiZJJY1NX
YvDwQ41FOIIpXBM/WVkmlcCfHLzfRBpE645SqfaHtKkfLLOgTt2SvMhAz+OsSJIZ4/25HNQScdN4m5aLMSJBTPWPtFtaDR4jJNiAk5lsHAPb6nEqJfFxun1uVVl++xcw
XQzPDspiGs2jpWF8nW680Fh5moeRLV3PGHwOEdxlgOO6+9x0TU1U+1qDZgR5SMheSW9NF6CKBuHLdrfZ8dEq9nYXqIPt2p0Pg8VUdhN0cpumMZoob2yeXCPcjJodlqG8
uv93rNO35wvvPI5Veojs0ESuqtFaC4ssy+ITOZpmGMdcJsaHeFu5n4hl8FP0qOuMddhPSfqcH8uV1C49OTK88Uq2qUlKZVFpnMWiTRCiuFsq/NG/OQFjdXnCdVe4ITZs
4NhFrwxGmyqHO+jR+TAV7fAXM1T58QqTeN91oiHyrYNp1Ad72tk28FV942WZ2xaeYQ262FdRbdZhAEPUCZR8cTWA9i9QCbPU5B59D5lvRA+jMkM1a1T4mqVsJJVRwDt4
2uZ3Ci/y+FaeQtmq7y7/+dWJAAmJf1z4Dx7U+CZu9cAEz7OH7NQB8S0bGD5jOdV7qfefUfdWnFSGoL7piGzzIwFfIWbye1EGKudLt+oc0z3STGeObs7fK9H/zE6InBQ5
VSHn0RFLrXTPvg8oVw9CKkkS5LmfqYehHudE0A1PFWLcndrloLewN4CGIZGy6NgEsM+sLOC3yGjoxPGgBo+9iSr80b85AWN1ecJ1V7ghNmzg2EWvDEabKoc76NH5MBXt
zNt3rGj9jD/aQjqEYE7O51XTlC8iCZEd/ZoeIRZe087dj57hhMwOPJmJyv4km1YfwOWJxWeuBRYMr1U4gNwcN2GAvi+fCvoALvwZTjluaDErxeMT3AL6h4ta8kIs97XN
ugpN6ETPpj4hVLqyDp2LJUlvTRegigbhy3a32fHRKvZ2F6iD7dqdD4PFVHYTdHKbmC5HEOY/sowCEiL27/l4o97YN+iWSI0zfA+1UPUf1bJVIefREUutdM++DyhXD0Iq
SRLkuZ+ph6Ee50TQDU8VYk0J6syb0HkrN+X9+7fDw6OE3gtIYGDNgDcBqq8eNgMjFRu9I0DRK0yUt0SF+495wP5lzTYULjYsWU60PhESCOXgSH2+PMsC5BIso2ErRJQ/
BFXSlXIeWFsYaMvHcrhw7d2PnuGEzA48mYnK/iSbVh/A5YnFZ64FFgyvVTiA3Bw3YYC+L58K+gAu/BlOOW5oMYhvchcQzVWNDRwM9L4dj+D+jMeCQKq1pYafiVJbi62A
BM+zh+zUAfEtGxg+YznVe6n3n1H3VpxUhqC+6Yhs8yPDVdVmVRbhJ3mNcF/m4Sfy6FytstiMAJS6OKxs4ss8SCo0kjYRofXmlqdnWqJ/5wkAI4ZoQBBRHtx+lGN4m0Mt
GlxL7HpTVog9WnQNDno5rps8e8iOIgREIkjUYfkE/nsq/NG/OQFjdXnCdVe4ITZs4NhFrwxGmyqHO+jR+TAV7b6+9Jm+TrJNJdsWmvoI3y5w5b9zLM0oGaBKUNCfao9H
tpKyfRf02/8tHqAq0NZuOtvqcSol8XG6fW5VWX77FzBdDM8OymIazaOlYXydbrzQoz/ttWCezdBZ7O90wmDmfgf8qXTAosUzPpYqBgl3UMTnIgz052WWswq9py7tYm8L
lND94lvC14gXu5leKvPbMq0ft89Zgad+KiopbJ3ocloKDLQ0qQCNovUuexI/JyB5KjSSNhGh9eaWp2daon/nCQAjhmhAEFEe3H6UY3ibQy1FJsbDk2Vubza87qqnQf3F
TJO2jrOfAJAEu8OA+wNJc12ZHHqmmtpAD/dRBL2J7QY4LQmSSAAfYL8ltwPMLaPBg3CVHoO501YobN/E5CPSgIKtsbiPCqssefp/yk4KOvRdjGzPzCt6lpGTxoB4ny+G
wOWJxWeuBRYMr1U4gNwcN2GAvi+fCvoALvwZTjluaDEc92IoaGuRv53jVjM/XPhy5MTHwCPNcns/aMRXjDbE3uciDPTnZZazCr2nLu1ibwuU0P3iW8LXiBe7mV4q89sy
dV+72ihfJW+e3HSNppyK/HEKFurvijIePthr7258jfkqNJI2EaH15panZ1qif+cJACOGaEAQUR7cfpRjeJtDLX+/OvGaGkWqdwFNiHu37WGuPFI+DVmUuL23nYlUsC0/
OgMV+x+76m5kxq6xL1rTZ+DYRa8MRpsqhzvo0fkwFe2q0NPcUFOMNnI0NuGrNPsSbnpoD2U1vqLsusnlUlwyy8oo2YfC5sH4iom1/1pAsmQ1gPYvUAmz1OQefQ+Zb0QP
lmoafi1Nfwgr4E4H3We5XzxVUuannxlAow0Y6meSL3TR5ShRIl94UvBsC1M5FJnJo1gqsdht9Ze0xE4OhuKcW5qPMxQfJHGlEqn2qRdUBJVYoW/Fszry4r0JGDFQPDXG
3A/PxgQYWgYJCytdn1VqUUSuqtFaC4ssy+ITOZpmGMdcJsaHeFu5n4hl8FP0qOuMayRhcTvR+d1Pbq0KdHU+ikdsTxHSMe8UaREA9s/I8YHsKeeaosEtPkTXFlIkXLOf
Y0mtqfRN2CloK4qBE4X/4cJ4aVU78MKCa/37RhMQ4hOhG5vJg5WA+fJ9sGgQv2HXG7pKpCz4AuDeEaRVp3QBot7YN+iWSI0zfA+1UPUf1bIHeKGobkNFyICQHjdr0EPD
WWCUWyq35NK7qqvL+O8qp5NbJBWcLYn7+U9/dE6sWBgB/bTut7KI4Tlh0MlT/S11FwkL2MtZisqd4/4zNjQQjM9zeakjjXO08YrecceHhPCiXc0NsGATCVp44IdbtV7e
Jz1MjxVV/HCqTvskm/mtyAd4oahuQ0XIgJAeN2vQQ8Pf2imKTfKRZ4eHbBnRNOXf+EHeVa81KZh9tvw1g+xMj2PEALUPFYF6jIxgInHejThp1Ad72tk28FV942WZ2xae
dLdtAEEnoTpjlAd52mcoxryxZyoSkPjOGWq6uY7CcYIoVHIKMbS+apsVZ6zCe/um7CnnmqLBLT5E1xZSJFyzn1SPwgTg3cdPSQS7MJl7J1ty/FYiAq0NXF+bfoMBsJb2
49PHyEUG9Gu9CseBL1Oq56epUfO+sm/kH+yASsCcF3jzlXAMOca1bzJisz/Tg/MnTPzLbu5v4geqQIr0eWm0NLSi42CibOM+/jEPGNo3WyNgAhrNvay0TTGuapxl7jOo
hjh6VuOXsNglkg04TNb9RJB/keYmgETpbFXygYEtO2rcD4apH2OU4kvJjUZnLJai3bElob40YEeoOIrZkJJTRD5oH5zCUnMAelN9lh1ZIOtmnyGWhoPgOZOcoCjnWlJo
3rdgMwHcs5xHKxXHDvdw0B+Wgwy17DJgNwYvTBm6LEgOiqkF9qUac4E5xwUkcdo13tg36JZIjTN8D7VQ9R/Vsl1R8yqDM078dDcdDR4Hs4jAXGeWmG8DVA5m6dL1HzeQ
5ZBiV3VB2X2hGAPZveyvqE8MDui5v3xtWO+Ab7T6cw/KKNmHwubB+IqJtf9aQLJkHzq5I6Ilq2y+ySKyzNq4nNk6Hv5BIlMNJ0kkQsNGnWoWw45NEUH2I5N3JHS+B3pb
3KpllSWEhO45sYm1KQSBa8YXFvVZKw/M73W+ltqjA24Ttrf84tfC85V7sqdG1yDWT1hi/48+omI5Iz5aXmCpUB6tKuqEDos1vDoKMegWEpKSHQiCdMpUhxUSWsFRcC9L
WBmclKMKWaRQlobaZUOn3MNuAjVtin98gHP2nwzaHLTRqlWISeXWE1ZKSa+6wI2rmzx7yI4iBEQiSNRh+QT+ezaiwLlplvjZ8o5ulL+lPWFZktvzHr5M1LwocIsQmD7A
I7OaTXYPtRLc4QusmiLfAbrSoXPPi8slp7PnhvL6SqmODgnxiXLheX1C76s4ubmKrzqys6hXw1zuIEwzpvo96HyHrJmgWGMcckTWLzR8Dj3cD8/GBBhaBgkLK12fVWpR
MKDACeSl9X6kjJe6jBqOBF/n8Ps9fl152CsOnK+aJW5HbE8R0jHvFGkRAPbPyPGBIHj0MFZ1pwX1ge7/raunt+C/tMk2zQPsZUbgHL1MkAoxYmf9TfvieZq4i1+4laBe
PpZsfBeM+mM9QXtpuP9NgJyWul+lrm+j7SaWdEqKSbVL4L2PBHfUHgQXHFerQY2MuY5z/UiHUqwsHvmOrlepRP5i+fvImwIiY5MfXPgdne0hGSFkulUckraU6giPzmJl
40q769Gv2Jj/Vz6OZRaALlbjsPeUkDv9UO3yj2H0C5yRMlp57brFf5LMWB0uYJwPww5AaTDDLgt2hMsUC/7iQDXRcL8e15Zs2WhMrBcQsKsH/Kl0wKLFMz6WKgYJd1DE
n8l5SSf48TKc4bTmBS74BWYs1XNv7ANxadjjWhu08mnVKZY8BnW6/zceu3wdu/UugBUXChQW4jk9V/40iULYjVvNAhueOdBJ4tOcLDU7Zb/GpHQlj5vBkTeSdkjOG/iS
3A/PxgQYWgYJCytdn1VqUTCgwAnkpfV+pIyXuowajgSk6sbNABl7K4hi8gQorKbXi5IpdFCcD+FVTbzsNb9+2aoTeKc3MfpwxlYlT8b2xwzvE2x9KdrA+nTjXyN2og9Y
cyX9ByKAb5LGOtrGlm2Ipxk2YQ3HQLPxuqXw8Ts+lmHZQldFGn1IUczOHITjQxQw/ljQisGm20MyY8foiR8+aI579XgaI7bLzpt/IOgkZQ/8+Saii5MakJYLxwpFxLYt
zvlkrhGs3RdsCM4G6GslFK9jo2vTh+VrXh9Rvp62ZalebJ+lz3gZ4J61woMiX9PpQAeMBSljlfAPAplTtMJjJht+KEDPu5URuDIIaTga4FzRIUb53MjMip6hQNhT1j6f
UQ3RcVVLuo8f8A/DJ0FOse+PdidNLzEPa8sPQvs0FjxIHqOfEHsLTpHSbi5HZyKyUZ8q+yz32SQAWUEBzAqfBni2ib5Ge8dax3ceRcrHwlmRJkmFGi/Nemccelu6M4Va
N66FNCoreQ7Y3+8bVYv0SJJ1XxYpJ4CBzJILILhMHsdAB4wFKWOV8A8CmVO0wmMmG34oQM+7lRG4MghpOBrgXMHWAZnZHZi966Wo6CNuUiDCeGlVO/DCgmv9+0YTEOIT
kTJaee26xX+SzFgdLmCcD6pS7/dxgvBOvDdq35b/C7Stlj5d1KQfiVjqiZJJY1NXfZvx/gnzd/NC5eryc6kAgUVXkdoO2Tahs0B8xUhC3CPr7YGHIrBw79ZVXMMfc9jP
mD/pBVcSn2m3rxnBQkkw0j2EirCi+wPmKXQovMUKZpEHGAWxAby5FbnNeZA5/rVOyogm0Sa9h4GMq195YwJtiEmqxVtUu8ZEDInZa4B5wo9m/64/Ch1sitprKBWwMqzB
knVfFikngIHMkgsguEwex70MlzPdZXYbxoHjOnskS+3pBPsLc+YXB1Nh77ougkYJh18/rZe+XKMTl+Ck8SldB5J1XxYpJ4CBzJILILhMHse9DJcz3WV2G8aB4zp7JEvt
6QT7C3PmFwdTYe+6LoJGCcMBUSLi3Sc6sR7Ti6N7EWeLyr6lAMTJ9WMf+Bi1PTyVYiHwckR7GFVhNv208iXw1+kE+wtz5hcHU2Hvui6CRglizBcAYtI+hrXGaLBh59uh
DT2KOrsT9gjx9wo9umnRP1HQv13R/YBLPROMHcAg1rJGHutkWgOuFpvQ/kfxDqH5qXghEQ7eaItwNKIaFBqiwK2WPl3UpB+JWOqJkkljU1d9m/H+CfN380Ll6vJzqQCB
VB6LcGAlTJg9UXiGkA9z5u3JSw4kPcJLzlrtLMiwITuYP+kFVxKfabevGcFCSTDSJW4b06ndW5fw1wk1VNps1iCM6sLGTrOHCPsGmwUvKtzNLBK42KSKL0/e7GM2D/ml
JbrMmTSyj9n+Q7wjTtehWoxLBfQTrASXbWueBcmb4PBWBg2q2AiZrAIew0p8jy1pjevdvMzufYvPTi4Rwxa1MiW6zJk0so/Z/kO8I07XoVqMSwX0E6wEl21rngXJm+Dw
K8JwWSHY/ZEURnIAGPwL9LF70n3BsRHmaaeIB1odgNVJqsVbVLvGRAyJ2WuAecKPFXYR6m2Z6aZ0ZwD+pL++3LtOvMO59rVDABk4dTMrZHbjUWd8J5mQUmZonBqVVrmE
SarFW1S7xkQMidlrgHnCjxV2EeptmemmdGcA/qS/vtw10XC/HteWbNloTKwXELCrsxUSRz4LeHjIB872UD015srdDmNmjSh9JoZAcQbwteTT/QlWbTbsaIHkcd/f7edx
N8/eWrwUT8o2kk5CTIOY2yaoh6yxFoLwHjXjWL1I4i29hX3tY7DdCBs0O0A8+JXS7xNsfSnawPp0418jdqIPWNUpljwGdbr/Nx67fB279S6AFRcKFBbiOT1X/jSJQtiN
IgQF4am1ESkUziUNq6miaSuOfv0DOXFsyHGNhLVXXYBHbE8R0jHvFGkRAPbPyPGB8gkJr9PNvv0l0V618wpLyzSxPFJzcVv4lAwB0CeOj8ldGpI9lD1MNItB6JWesRpt
R2xPEdIx7xRpEQD2z8jxgfIJCa/Tzb79JdFetfMKS8s0sTxSc3Fb+JQMAdAnjo/J/etVm1E3LyYo7rRPANAXj0dsTxHSMe8UaREA9s/I8YHyCQmv082+/SXRXrXzCkvL
NLE8UnNxW/iUDAHQJ46PyamptbmsfNEs8jaA56aQpPVPij7JwWM0tqL57l8VlYPPPBtm2eOc2T9zCe1AyEO6/G0xohjSzRs8thLEX+w+oH+2BLuVVekb0Xyl9Itst/a7
cyX9ByKAb5LGOtrGlm2Ip3zGVGSJWJbJxSnCM1PEoA3Id9f3QS274L9HFZKZo9DyxnSX4b1Qcva0o662GMby64CmNxzirTYd7fXcs4sXVISE3gtIYGDNgDcBqq8eNgMj
H5TDSK7OpRLyCv4fddzsex7SS2uCwgZP0KSay+QnUSGN1lLHmEziY55ufOqahEJMNdFwvx7XlmzZaEysFxCwqyWIL4I9xEJWIo3aet415yX+0T2IRNcSxDgxcor2opWG
Rpj/0IKCZOn8728fCke7+2UvXig1hiXyhDj94sIVZvg1rkJgx2snt/UF/MNYFEAYVCNQEFtzTjQw21nI2NiQQjpFaV9ZjyW0vKCFXl3gH29egkbmb67G8/zKxK9/bVCb
4/25HNQScdN4m5aLMSJBTDCh2BroRwyuWmqQZaa5pLY6RWlfWY8ltLyghV5d4B9vrPG6GLH/hjh6dRqziORoshcJC9jLWYrKneP+MzY0EIwXqP3PaPaURtHGf6ttI6ja
AuocZcRiEJ9sgcbvLV3atv1zFW7cdgpnZDL2wZ2XcCR/FwudDKXKnFmdEuYD3eGwCKoKmtxpiX6tKsVc0GpoSh7SS2uCwgZP0KSay+QnUSEMLu/zS/sOcMsa8cz2ZsNy
sM+sLOC3yGjoxPGgBo+9ibRsbNjWRvUmvtFNZE17xy5d383aHFG8pLoRz/CmKgF1mERD6Tgr5E5hZT3u6IKxs5s8e8iOIgREIkjUYfkE/nu0bGzY1kb1Jr7RTWRNe8cu
Xd/N2hxRvKS6Ec/wpioBdY9PzlpLPjpIuaPfEQo6uRWtlj5d1KQfiVjqiZJJY1NXCe/ZROonP1e6KAq1WDD52gi9JRYLPs8uhpFWo8kbyAJfU6VO+iCXW5jm+8B8kGmv
rZY+XdSkH4lY6omSSWNTVwnv2UTqJz9XuigKtVgw+doIvSUWCz7PLoaRVqPJG8gCdV+72ihfJW+e3HSNppyK/FbjsPeUkDv9UO3yj2H0C5w8G2bZ45zZP3MJ7UDIQ7r8
bTGiGNLNGzy2EsRf7D6gf446BwW7AaEpqAwqUsdfPFzNF01DOloU4IgZ7d8HzUS5c3dmzCJOcvm+4QBVQ18Y2gswNYIgE/X4ilJCL7Szsaofn4Rnr93kNGReh06LRfdE
4Gt/JLYNXcKFu4a8OaBRVMh31/dBLbvgv0cVkpmj0PILEltCxBmX0+vYC2xxr1Lu23iajBCwgP/c5j++AtTIa1QjUBBbc040MNtZyNjYkEI6RWlfWY8ltLyghV5d4B9v
yNyKVC1RnAxj6ja9iFmu6g8kxWRPpKAatSVRsRjAsz9mTdjTi7Eolx4cogn5X0ZXu0A7EV1bdj0SoV9IymjICDvEoqEeQfxkg5zPLL4ScVqQ3U9q3FAufoBEPwYYR/v1
evL3bvI4DtOB508+Y/7iNUAs+KqMWrEidEanZMnBPkA0GVfRPQVvXY1UrNzc1eCKYcoSV7/chJy3XyIdtTH3rDHeQyUVwiYqY8nauQP2mnB5W8Db7d5UBvCzdVCaMoO6
U7G5da5OCaYXvknkNwDKgFwmh57XKMvDFj89en4e4tJkagK6sB1dV5F5bp24LBYei5IpdFCcD+FVTbzsNb9+2YrbUbxq1zsLwzQKp68H+SlXWh7kS7mv97WX3yWLXj0F
x/TvyXusflafz5M7XP2cviWIL4I9xEJWIo3aet415yUKUTqwmEUCveNrHDvR6ahiZizVc2/sA3Fp2ONaG7TyaTxpw3c+8mQYZWRGe/aKJhXkADrfFuZyp8+RDkMIp58J
jwCqN4OYZvEfVGkCqweDt9dPiiF7BWEzhum9GrrdmrdPFZBOUjULwGNTIofMGhniouT0kb9746EvKNjS8ePEH90ERJysncLlt5pAkNIJoOwO3+nYmei3D6286yNXY+E9
YeGAD78OIzQM8DvTFZ+RReGdb/T/UfYaluo6tElKv9SA6zdkyg1WLuvKQUXMryF44/25HNQScdN4m5aLMSJBTGHKEle/3ISct18iHbUx96w6KBFQMXrKRXNBZJfVYicx
kOoC/wtscouWuE1hL3U6XanCkVaC+VIOu9QtB6Sl2YG2lI06FVws7R/e0mm0UfEWZEkljiuTsidH93CjhXspEDFiZ/1N++J5mriLX7iVoF6fk9ENsGC3nDK1Ftnfm1aD
T3uOYf81ndVatzKlsfwFeeNKu+vRr9iY/1c+jmUWgC5W47D3lJA7/VDt8o9h9AucXFt0jqoKcINeVahj1zU7b9P9CVZtNuxogeRx39/t53Hs5Fyl4GDxLVwW8EdmyiGc
69AvDo6xV8NUzYXGVumiuPqEzQZwm4zRhJz3DndtCS7MZllzCqTY6yz+HPMIFTIoAlHqFjm3ENdwQsx67B2Nr/fiTczBhFnVEmWnHxL4sfORJkmFGi/Nemccelu6M4Va
2/kCIcUfW+/KLSRTCF06Y7DPrCzgt8ho6MTxoAaPvYnjo7fzaC/Z9MtMi8MMs/4lG34oQM+7lRG4MghpOBrgXPn4dou/LVt8hGYonspLjRAQq1EaSO+ZWwV7cRUhbgF6
+oTNBnCbjNGEnPcOd20JLlk6ofNhz0GeBRaUDKdlD1Z9zSm8p9XzuJIfkz+RPTe54Gt/JLYNXcKFu4a8OaBRVHCBE8N//Qwi3gi6RXn1tFQBFrVPPqZPd4+4JZzI4Fv5
U9IkDqnzU3Au+xtSXEy79JM0VdzAHy0PshMtyrlZGEEqQdNgtnd4VWBHoVyrxvysnYIoIqJcsy9SRs0EJvehs8Fy30H41D4NqMkRF6n8CW3e2DfolkiNM3wPtVD1H9Wy
O9rl8BsN7e4CF/4e5Xs2uGj8ewgqg9dlJQPyPPXvxdYMw2Wi494QEgYtGUE2LFrM1u+ogQQ9aHf+oHmSxAELNTFiZ/1N++J5mriLX7iVoF5zgKTYNvm1fIUQtaYsDZFv
gFBKtWt1Txj2XkTqzIbk8rOtDqt20gCMNo1wHFOevZVdMVa3isAWX44lvJZB7woM9t/UjK2AtEi/+WlVoupiah9XgbOiqB9chVJY0lSJdNbKhutP56KtseqsBQIPMSVz
IcsIPWnSZnuVsm6Mtakl4GLMFwBi0j6GtcZosGHn26GBIRQGKEmnt9CNoBbHPULyklYHS5SBDoDTfBwg3BzJ1WUvXig1hiXyhDj94sIVZvg1rkJgx2snt/UF/MNYFEAY
WpuMDhdD8NerFopk2Zn7UwFGZjN5LwdFX8/rAk6mfC+AB1e3CoO2uQxxNQuHfg4UPhon2Ja6+717EogPQJZ7Clwmh57XKMvDFj89en4e4tLM8OSBu+ytQ/KWq8VW8skB
3tg36JZIjTN8D7VQ9R/VsshyniwebmgobwMBj/uMDfH6rNttf/2pI2Brg/C/kWoguY5z/UiHUqwsHvmOrlepRB/aSn+QfawrPSpZl56l7N8hGSFkulUckraU6giPzmJl
zgdcXjPmF9DaM+BGoM11L0+KPsnBYzS2ovnuXxWVg8+ngxsJXtbxSWJbn9fwoQEpww5AaTDDLgt2hMsUC/7iQB9XgbOiqB9chVJY0lSJdNbKhutP56KtseqsBQIPMSVz
L75jQ28u99G6gzXWp6w1Z1daHuRLua/3tZffJYtePQVyMLXJsQur3Sru1eD9gce1sQXd4sLWugduIZKjYlVRlI8AqjeDmGbxH1RpAqsHg7dhFvMjZAIYRjUP6qbaWioJ
LVzyL0eTV5i8SMk7EIMRRJ6XGw3Yjp5BSq6g1tdglMaRJkmFGi/Nemccelu6M4Va10ggbg5WinIhLK1axu5Hdj4aJ9iWuvu9exKID0CWewpbzQIbnjnQSeLTnCw1O2W/
lKPloq5LGBaG+UU3SRTQwIEo9/W7TJsV79ozl2OARJxR+IM9yscSquxGpxEeYS16sqy3gzfS/Ab7LSu1771xb73N6eugI9QosBXhV4l4rH7zpAg8diJ1zWjtUQM3I1XE
tpSNOhVcLO0f3tJptFHxFoCmNxzirTYd7fXcs4sXVITSLXwZiBQBSDcJYITFBioWJ8jd2usOekD7q+J8zf1AA097jmH/NZ3VWrcypbH8BXnPAv2gQzmbJvJ21upI04GI
TvbyRR5nuyKf2hYshUW+U1zFnvQRo8peIvmLqpfEer6MSwX0E6wEl21rngXJm+DwaBRKWnTzIEaGy9yO+1VgWjqGyANhyvX046ZIki3DkN9t3WE729ZK+LYBKpHOlbHk
OTl5MsSDYY2mE1Qj6KVvbw8mf3oXGvuu3tmstxsoT9HDm3dspN6QhgZcRoHZYSqdOigRUDF6ykVzQWSX1WInMdgabU6Op2o3VPgkmuZ1A9sNPYo6uxP2CPH3Cj26adE/
XMWe9BGjyl4i+Yuql8R6voxLBfQTrASXbWueBcmb4PA7h6AUKSU3+19pajJRvCbJyogm0Sa9h4GMq195YwJtiC++Y0NvLvfRuoM11qesNWfRZDB22KF8NGSOXY5Dh/mD
wnhpVTvwwoJr/ftGExDiE3ZDVV78Ye8EAdmLav5oWM/INwe3r226U0othOlXR6gNKkHTYLZ3eFVgR6Fcq8b8rBpLdeYknugJDJ429tztYsRfPJqP8tLqxEm6aXUzsXEw
7clLDiQ9wkvOWu0syLAhO3bSUdRyeugfF8jfyLD1rnWOh4/Jm52dgiX5lVBc59Ssd2s0Fq1+5M7yt7nnWhtBJKLmbbnTFBvmrPsKTM4kkD4omHUe8qWxrDh37ZiK5W24
11cAtaAO9BXMvrMB9ZhZlbOtDqt20gCMNo1wHFOevZVe7b1jtGUO4wCOVyADujKTff6nrtmOuw7XBBv8jcv81ZCJ5JE+YPF02xH1LbNuUCqxjR+9tI3HT4wmp82OanBJ
ydkFDOGgHPGptEROCsC9HOCuT3CqMLhvoWeyLn8TCmlhsWwLXHAoNbyYilpKhZNlknVfFikngIHMkgsguEwexwRrZyNQ490sUIcypjRTfsJJYNU8ifkn1umKEgDAuXoq
qXghEQ7eaItwNKIaFBqiwK2WPl3UpB+JWOqJkkljU1cBsfVDkycbYPz35xXwuJCYjT8dDvCSpB8LvKXHEVNtGXc2EUmKaxFqwQAYeiKQNUf8Q+EL/rFEn+DYI9fZMjjJ
VCfOSE2+lzvwL6JTgFtWmDxVUuannxlAow0Y6meSL3Re7b1jtGUO4wCOVyADujKT7kaM9Wyr4TMdNryQL3jT8Ge0KmmL/S48dP2BLR9cPkW5prDtMVhiHfJELcocL5ad
Ty5E2CINky6Lfqya1qiAdJr0Oy4Ve1uAgriGBBWw589TYyTerXB0su1jYcSlJ9giRzTtJyAvYfWbvtmy0g3mBG5Zc2C1aP4KbypRQQHrKLvrTKtOh9U4y4beXumFbqNv
CvAIiiNvZswqVu4wA7r4sOzzOnG81fWaUX2+9m5kxvejOl3OrqIimr/pWL01T2FCeOoVxWItOiNVRpo7nUfc5mc4pa72nWUGQh7HH2zGPRgLLFLaTFxY73WsApJEEiuF
VXqqn1B3lMst6anUmjV4Cfb/U/ordXxV6/vsKuSDm+OaR6J5ezJ0bgSSuA5M0y8R5o2GRkz6ceXx5Ax9dmnkxlTu6onrsuJ+KChkVI4ceh7T/QlWbTbsaIHkcd/f7edx
N8/eWrwUT8o2kk5CTIOY28jI+jBoeUxIqVHg0n3dBlLBztzsXHx/6zlnsdr4LC5n84/ivEzHZIw5w1PbgmdQlS1c8i9Hk1eYvEjJOxCDEUSelxsN2I6eQUquoNbXYJTG
7kaM9Wyr4TMdNryQL3jT8FEssSGm7ex9Or4nRj4+i43Zu/KeLpAl9F2UYWgwjuHy/B5QhOdW8YcjHbRZpmJqY2IGN0IkfcrL2dNTaCW8951PDA7oub98bVjvgG+0+nMP
1ac1soZgVWyG90sfui+canGgEgMQK3tqHmt8hD0eIXtoChyUa6ePsWISc002tmqP3tg36JZIjTN8D7VQ9R/VspsAFcYvXeJ5AydeL4wh6MehF/4pyJ1G587YJgMr7JlD
23iajBCwgP/c5j++AtTIa17E3k0Xh9M7lga65gUzMAOU3JRIWQHkgYdGP8ybClm7tgS7lVXpG9F8pfSLbLf2u3Ml/QcigG+SxjraxpZtiKcTr7fBIMYTkjBP05A0/fdG
kflnpNqaiUjqkgudb74TPZ8cYdZelJOjvPRmgkiwPTRWBg2q2AiZrAIew0p8jy1piDykPge2eUW3RxMBbR8zBvweUITnVvGHIx20WaZiamPxRJ4UvN7lyBOYsMY0Wyky
mkeieXsydG4EkrgOTNMvEYuSKXRQnA/hVU287DW/ftkb7MHSyef2akVwMUiozokOVjBx8Q7LdGHA00iZtWKT06l4IREO3miLcDSiGhQaosCtlj5d1KQfiVjqiZJJY1NX
pFvdKhe0HrrxUjWSj1Jb3jj7CeshxG7njJ/uwUq48THGpHQlj5vBkTeSdkjOG/iS2bvyni6QJfRdlGFoMI7h8vweUITnVvGHIx20WaZiamP1tk9ddRmKd264qZennDWL
23iajBCwgP/c5j++AtTIa17E3k0Xh9M7lga65gUzMAOU3JRIWQHkgYdGP8ybClm7SiE0m02CcNUR78L0trBVRMf078l7rH5Wn8+TO1z9nL6uYdsrO1Si8zCZVFrqFfgb
BDhwGElGa586AhAnir2bRjdajrskJj5gigfPotoTGm+cOMbBvWZ+5UXESEsYnHnakyjNbvtloOMTsWlhkUC+Si0L/PBcnwItEG4UuvXgSfiH4t+whMz3dhup05fk+MMa
ZOPBketMLMQJFkuna2gtQfoiFHqHLUjtUhhvqeAmOo0wZfOBL6RwkW466o/J2HmIlNyUSFkB5IGHRj/MmwpZu0ohNJtNgnDVEe/C9LawVUSAYoD8TO41bl+w6pbKnASz
yQgzuZRYFx2Bu8ZGVHTzHwQ4cBhJRmufOgIQJ4q9m0Y3Wo67JCY+YIoHz6LaExpvPxk1OiO1vwOjY5w940pnByc9TI8VVfxwqk77JJv5rcibABXGL13ieQMnXi+MIejH
cGR4YExAy2v3hbu5mfwmxHLD61xHv+ffRNZQxfXwHjO5jnP9SIdSrCwe+Y6uV6lEpFvdKhe0HrrxUjWSj1Jb3jj7CeshxG7njJ/uwUq48TGgb5NCX0h2/ImG4tzBlm2A
Y4RvCbYmY68ETsPzFuDUL5TYV8WLI/t956zxFyTZyjhImzE0t7W06yA/+OvXsfALpwGYnuSXVW207/6RJUv2EJDdT2rcUC5+gEQ/BhhH+/UJRoqfMVUhlqF/ygAV7TW6
1KCfAGTUW9x2ns+0dtT1r4uzYLgMEED2ij4G8pG0slHKiCbRJr2HgYyrX3ljAm2IG+zB0snn9mpFcDFIqM6JDm3OgYGKzLAsbg1nUa8XFnuQ6gL/C2xyi5a4TWEvdTpd
FPrtoEKuaoOHL4SYffSTp0ibMTS3tbTrID/469ex8AsLcjJsZquSzdnnNfvuIDin7uaCuyDtKa0z7wx5n6LJ+AtXUTG2LpkqYrGGVPp4ov/8HlCE51bxhyMdtFmmYmpj
H1VqUNIfXhE0JXsgEQKGsBq+EfAZ7a6D25O5Iqgs7DYLLFLaTFxY73WsApJEEiuFPEMVzCrv61pC2Vt0VppDOC8Lvy41m/VnxgzAaRIGVl2Kq59VLpM5SEI2mM4luCdO
TE2LdOmo2nE974iJyIl7kv5420q7PC5ThgpLq1L38u5ImzE0t7W06yA/+OvXsfALC3IybGarks3Z5zX77iA4p2gUSlp08yBGhsvcjvtVYFqIPKQ+B7Z5RbdHEwFtHzMG
/B5QhOdW8YcjHbRZpmJqYx9ValDSH14RNCV7IBEChrAZTKFPPuzuYKhtRkZk1umCCgy0NKkAjaL1LnsSPycgecxlw6pA73AIxb78JHDw/qtv90RRDf67G3YUVjVlvZ3B
N66FNCoreQ7Y3+8bVYv0SJJ1XxYpJ4CBzJILILhMHsfAfUBZw/m1qzBb7TGapWC+1KCfAGTUW9x2ns+0dtT1r/OP4rxMx2SMOcNT24JnUJUtXPIvR5NXmLxIyTsQgxFE
/2+oX+5uOUAm4pnqeyknWAnvLZzqPbE0VxYuuo4ZtxxHFpOt3I8Du+3l6G+SyyZdKkHTYLZ3eFVgR6Fcq8b8rDeWEXXDgUAgj9Brh/+athcHzeD5fVv/bQxZq07acXvJ
T4knUM/Lhz2gEK3KmIzVn97YN+iWSI0zfA+1UPUf1bKbABXGL13ieQMnXi+MIejHZUqEbINdVit7b1A0i46J6zxVUuannxlAow0Y6meSL3R/RVStluUJobBTcM7zgJJi
Ce8tnOo9sTRXFi66jhm3HHIV/EFXjdN2whqssl5hpZT3h/qIlGioZWR7wiqSzzvIi5IpdFCcD+FVTbzsNb9+2RvswdLJ5/ZqRXAxSKjOiQ5ci3N/QYM/ULNS4liqYrsK
wwFRIuLdJzqxHtOLo3sRZ4vKvqUAxMn1Yx/4GLU9PJXAehyYd2DpEeB4oLcEswZ8HsntpYqWgjYCbOKHloIS00tthOIIO3yJR+oDaBaCdDI+EVjclhk5GMVNqGoHM7qC
lLO1O6RNTMlG7Us3l1E63wnvLZzqPbE0VxYuuo4ZtxxyFfxBV43TdsIarLJeYaWUu068w7n2tUMAGTh1MytkdsqG60/noq2x6qwFAg8xJXMb7MHSyef2akVwMUiozokO
XItzf0GDP1CzUuJYqmK7CmLMFwBi0j6GtcZosGHn26FC2SZ8RS0ftOftsC5mfZf7LQv88FyfAi0QbhS69eBJ+BhbW5Qoogyfi4zw6rajWKy02QTVdvHB2XpEHJ7t08qr
MWJn/U374nmauItfuJWgXk/1dxZfsdKzNAj1vlm4FucHzeD5fVv/bQxZq07acXvJ/59nCH7jzBbGnCozgXovCn3NKbyn1fO4kh+TP5E9N7mALFP3rF4vLbSjTQHuSXxR
kflnpNqaiUjqkgudb74TPV2oldFkMcaEDzMQL8ixM+kPJMVkT6SgGrUlUbEYwLM/JQIN6+P0OMns8Doq3JiZIGuDqpaWqGgn7N535YjaGkvNQp+wHBorpK+5DyVo3fET
wnhpVTvwwoJr/ftGExDiE8xlw6pA73AIxb78JHDw/qujbf4MF/0/CXFqlQRluXZWZzw8SoLjjdgHnAey4TmTOROvt8EgxhOSME/TkDT990aR+Wek2pqJSOqSC51vvhM9
lWrr1vBFJLFh5+31QK58N48YemkG3G0bemgoHEEJmfLSTGeObs7fK9H/zE6InBQ5mwAVxi9d4nkDJ14vjCHox1NMnJj2pRBpyHAkYpQjqp6Apjcc4q02He313LOLF1SE
hN4LSGBgzYA3AaqvHjYDI+ndD52qJevDBVizUspGz7oHzeD5fVv/bQxZq07acXvJSaBiTWbTYYrTqIhF8+bTGZFca0DiazmbKzbX2pIzjhmYY8E6xge6LRDm0SgoPK8Y
kflnpNqaiUjqkgudb74TPZVq69bwRSSxYeft9UCufDfRIUb53MjMip6hQNhT1j6fUQ3RcVVLuo8f8A/DJ0FOsZsAFcYvXeJ5AydeL4wh6MdTTJyY9qUQachwJGKUI6qe
x+3FlrY6oxwtmNL08m03e2gjPa9L81g3aFJI8x56i+mkW90qF7QeuvFSNZKPUlveyJfLoc89PHHBPt6rH1j7f/6lDkKM06uwSI0qPfh+/4zAa8LG1RH5K6YLHhV04v4y
z5Vr70Gi0e2SnnUQU+Dsr2uDqpaWqGgn7N535YjaGktSMwgq1rkzRDOh/H3oVQEI1SmWPAZ1uv83Hrt8Hbv1LhKEqu5eY4moQkLgYLOWYjLQ/sOUNcTkGa/HJWED3bdx
/uxsToGU7DakaHEcS1GqTE8MDui5v3xtWO+Ab7T6cw9tzyRt/QcIeoko81IrEZC+nRTm8mCn2/d0gcjbGJ7S20D0W+RonFDLtX/JqDC0uwTqCVH7mTDDRcUq7S2j+cYO
sboBP/MOvcANSggSltIArPBvCU5m17s27y6hMkccqJXKiCbRJr2HgYyrX3ljAm2IgjL61U8H5kSH+Oyq/GhmLB+C3GLxPi8ZoYk9h60oIFF3mdvpTRyo9LtrOcui9Lfp
KM0/KjiZFfe7z3jASnt48sThYsSTfayWwVBKwC1G13oEVdKVch5YWxhoy8dyuHDtIr2mVvCq+iJ88Tfbqs9B90wa5kxf67wTtES6rinjigK1+uiJ2QafNeTiimOstzYZ
KUBpdcA/ZPpqHuGhc1yHNbG6AT/zDr3ADUoIEpbSAKyqicTn295ufn1WI3bLUkzO3tg36JZIjTN8D7VQ9R/VsmaOHwTW2N3QQsWXcrFqKAnnIT3Mp5RaJoYrpLXSRAlf
i8q+pQDEyfVjH/gYtT08lV0JzgHrSisTNI4lNrro1Bh4CgKCLqsqkXPFK2pw9ClNDyZ/ehca+67e2ay3GyhP0aJmpuZS0gFUxHjGcaEa0xf3I6QEgtdqrEC8yahx268V
PWSC7M8w31wGGEaPXd72mPcUdu8ffv1BRfuVhcaXiUqeZevuxuQ0heAHucWv+L4i93xYpbUg3++BMcj2bnPATvvK6UoFI6JENGSIFUP2fJKYdEXXd7Xu4eLXFj1Rz70B
xvbRFVL3Zsn2CxcQTilwHVxBjZ1YR2iJT0kzuj6ib3PCFyStaJp4ZS8JXNzc6kLPrpFbU7jx3lJiX5lP9IPEQsAEeTn8Um5ebkClyOxTWbpMvyT+sGvO46YMnHtQGBBG
Rtkv5oPUN0pWdD3TY2HL9fnVDFMoyssGteq4IV4c3SzEHIdud8oMs+UqTLgX5JgsSASi3YQDqHhYMur2b0/W53BFbG5YOM22Uqd/rK7SSLJnnN3kDz5uD2mGg+jRx7Uw
7VgWGw1E4gRpJwUmLvyU2Kt2ZCl1ztiihVF6gSdAlx5RQ3Dk70dIJMD9tmqpBYl4clCjkxpDOzajk8W4JmT/DylAaXXAP2T6ah7hoXNchzXJ7OQw929ijH8IssWq7utl
PXHMYlw3k9AGhFIDJwtKOerWeb58Xut3tyAiW82Nct97xqCUNVolHb1aY0m/p4+L/yGOXXDdEmQNj71GofJkkbCu/eO+S21XWnhmPN8uxtUucE8tsKM4t/lbjxbOt2VH
JEGBnRHtY9akbcmpB4BCTJfax4KzqbhAoinP+Ix2Y6okH1IHf65Ew/TrlyLgdaMLJU6U+N5TpzlISBg7MYyphE+KPsnBYzS2ovnuXxWVg88kH1IHf65Ew/TrlyLgdaML
VvnGVjDk79i/tgh33rCIrt7YN+iWSI0zfA+1UPUf1bKNhfhcuO6fbCHdKxfnvGTzGtCt1RVgh0GklKucVBg1SEdsTxHSMe8UaREA9s/I8YHhB86IgxbRdF4NNcusea7x
78fLXly/w7CQgzlGwUOefgssUtpMXFjvdawCkkQSK4Wmxrdc9nBI97K7fCFNCdC6kyXT7dDzYI2x6qIhDdmFq5DdT2rcUC5+gEQ/BhhH+/XRruXT0sePzV7TTEDVF9om
h4PZG9YTnRnmCLToaS+kLoTeC0hgYM2ANwGqrx42AyPLMJKOMtEdsQB8f+vh1wovCYiA3SWhG+wmVk25FWvAnfd8WKW1IN/vgTHI9m5zwE77yulKBSOiRDRkiBVD9nyS
0xJE4TmwPwOLW3RyfvdwVcQ3pjbeT3oHeYQWIJn5W7Ci4EbubW50Tt+cDV7ASNMLeGy96KZtr7zJxHgom9++OaHmbs763+meI6ndZNl8/LcejLrHZJrCotJ5psNKy0Ua
eGy96KZtr7zJxHgom9++OX7e7u+HMO6QvQK6STAUkklwRWxuWDjNtlKnf6yu0kiyu2fijNHoSmv0fF8tcFgwPIhk01eXZxuY0toMAhkBWJgpQGl1wD9k+moe4aFzXIc1
hoZlICPJIv6ZsTXmOWnFgKbJGcgfKq78G/EyH5Uvvbjq1nm+fF7rd7cgIlvNjXLfe8aglDVaJR29WmNJv6ePi6ZDWdGFme1QnbY8wwjjoTqwrv3jvkttV1p4ZjzfLsbV
LnBPLbCjOLf5W48WzrdlRxOCN9FaKVWdjvS5yzR18+kPDjssEpVuHSpP2AAlY/f5HPuhzJZjrEEFDaNRawo/tBuNXJ3FRZhIkeGFf0PJt/vKiCbRJr2HgYyrX3ljAm2I
hc4jSwzDsq2W8fvr8FGgKkp3W67k0JlWxk4IKjhe0W31p78L3zb9NpqeLEVMWduFpsa3XPZwSPeyu3whTQnQunWt2xVyPWUqSZN3xLI/Uqq5jnP9SIdSrCwe+Y6uV6lE
kG5pe6NmfLEfvLd1MVathsq+sH18wk4c3acIfB1hXLJHbE8R0jHvFGkRAPbPyPGB4QfOiIMW0XReDTXLrHmu8dT78l2HWDe9cuEzitIsILmQ3U9q3FAufoBEPwYYR/v1
0a7l09LHj81e00xA1RfaJp5VNX/o4qJ/u4T7d05W44yE3gtIYGDNgDcBqq8eNgMjyzCSjjLRHbEAfH/r4dcKL6V5J2+YWrXo8/YnB9OfYIH3fFiltSDf74ExyPZuc8BO
+8rpSgUjokQ0ZIgVQ/Z8ks3CBBiUr+I6u+e75FKXQt09ZILszzDfXAYYRo9d3vaY9xR27x9+/UFF+5WFxpeJSkzKF+Aui3QeOz2vFWzCBG4PJn96Fxr7rt7ZrLcbKE/R
omam5lLSAVTEeMZxoRrTF5inAFbljrJ8gobYk/SO1SiungKTcA6QV4Is/cpALFjriBmMN6NOhA6tWkKYT/hdjXvGoJQ1WiUdvVpjSb+nj4uwtZ6Mpj0h9I71+kGQcMZq
8ihQrzc9RAf0qdUSS9yBq3vGoJQ1WiUdvVpjSb+nj4s+SMFSqKvGdf2cDM1W6wBRKUBpdcA/ZPpqHuGhc1yHNdX/xBbsQD/jjPOZLi8VNQpFQyZGjCAoxI91wN5yI/CI
sK79475LbVdaeGY83y7G1S5wTy2wozi3+VuPFs63ZUfj/kGWCeFn+3/reAeHGf4FDw47LBKVbh0qT9gAJWP3+Rz7ocyWY6xBBQ2jUWsKP7TwHZMk94mhkiC5FtMu+hMn
yogm0Sa9h4GMq195YwJtiIXOI0sMw7KtlvH76/BRoCpMgF4dNwiw9iaAkdz0P1vNUQ3RcVVLuo8f8A/DJ0FOsY2F+Fy47p9sId0rF+e8ZPMY5+3XaT7B1b1XD+LV8Cbt
wnhpVTvwwoJr/ftGExDiEyQfUgd/rkTD9OuXIuB1owvksAGo3c6pLovIBg+ZvaNlko6BC0DmSPNQL26NcLqr9sswko4y0R2xAHx/6+HXCi8KPj6LG31B5Ng64j4jV2fx
MWJn/U374nmauItfuJWgXnQCzDTe0oYwJ8h9T55HNTsa3nKn1m1eAs6acGz3e4OQkN1PatxQLn6ARD8GGEf79dGu5dPSx4/NXtNMQNUX2iYwLmzBXg5M9/1lLiQG1ktl
BXHrW7Oo/J3hRT6snWR9NPvK6UoFI6JENGSIFUP2fJKBPi1c6vo1t52SfL66p2z6FQo0mTEQFMdX5ZzLD+847vcUdu8ffv1BRfuVhcaXiUq0e/SmpSCDWWexT0vSiPHw
DyZ/ehca+67e2ay3GyhP0aJmpuZS0gFUxHjGcaEa0xeX4p6nUiPVLpcltfNH3Dv36+2BhyKwcO/WVVzDH3PYzyeSBRk8Qoa9QZhpwjaZVzFnb5go9RqQ1BlHQvV302Xt
oOe+sYVgUe6KpWaZdisLy93kMlt2hpuwmrL2Iuec5CEWMQV4pFeNi5jw6adR5JqaHT8A7mj8quFIny/IsvpgNnjUaTs4bNZSDZx49JYuOgAc+6HMlmOsQQUNo1FrCj+0
ZROfPQuPEbivihWSxVT8DRCrURpI75lbBXtxFSFuAXoc+6HMlmOsQQUNo1FrCj+0HVgNRnKSc89h1dvJ/Qun47Cu/eO+S21XWnhmPN8uxtUucE8tsKM4t/lbjxbOt2VH
6X8FMMM8DKX8sHMwUZVWcsqIJtEmvYeBjKtfeWMCbYiFziNLDMOyrZbx++vwUaAqqcZmPhQSrswLa1/EtTIrq1EN0XFVS7qPH/APwydBTrGNhfhcuO6fbCHdKxfnvGTz
KbqDJjHyeykTvpqrFtm06MJ4aVU78MKCa/37RhMQ4hMkH1IHf65Ew/TrlyLgdaMLTuyZrUS9IuTQ1/ZV+AnbgJMozW77ZaDjE7FpYZFAvkrhB86IgxbRdF4NNcusea7x
JsZRKOL8VcSSGgx2J4x1t62WPl3UpB+JWOqJkkljU1eQbml7o2Z8sR+8t3UxVq2Gd/aIcO6A7I92tH7hjh6IlEcV71y+w1MoBsGr42/xUojdkQWG/+pskdzIE65wuQHC
Lj0q/w2xtMeiaWU73+o5ahcJC9jLWYrKneP+MzY0EIx6DbwgYg5GfZdNn/asjxtwLTSs6Y0Oo8pAqfRW9LrAcZIc9KIp+IdTN6r26o9igSL7yulKBSOiRDRkiBVD9nyS
UJFEeMxd1TGhUvWrfTs0dZeQ8U+1pQoV2yPWTHfMvHWiZqbmUtIBVMR4xnGhGtMXZRRgRAy5QhYGcSNgWOauqvbeshtcbJO9GascshhESO8nkgUZPEKGvUGYacI2mVcx
637UUiIX+efGoTlwPUnY0b00aaRly14jkuHe525h4Ojd5DJbdoabsJqy9iLnnOQhOZY6UWSU0dm3vAANZca6K0D0W+RonFDLtX/JqDC0uwTqCVH7mTDDRcUq7S2j+cYO
lxzyzLsRn7inGC1uaX/cm5yB+APQjLlz7V1eSSP811SKrMHJ3VgevogEJrXuKyN3e8aglDVaJR29WmNJv6ePi8DuRAp4Bujfo1/HoA1svrkNKIS5/6HJvZISH2E93wdK
jYX4XLjun2wh3SsX57xk84mIBRZR0VRGv56/INnf8rXSTGeObs7fK9H/zE6InBQ5jYX4XLjun2wh3SsX57xk8+9egci/x5/1D3PNY/YN6nXKiCbRJr2HgYyrX3ljAm2I
hc4jSwzDsq2W8fvr8FGgKgYvigITRUNAqS2uNX3WSWHCeGlVO/DCgmv9+0YTEOITJB9SB3+uRMP065ci4HWjCxPMyz+QsxAEKf/J+m9xFtmTKM1u+2Wg4xOxaWGRQL5K
4QfOiIMW0XReDTXLrHmu8fRoTwUV4qO88/DrDlYApmKtlj5d1KQfiVjqiZJJY1NXkG5pe6NmfLEfvLd1MVathpNZManapWwMvqu9CYsSgDKLyr6lAMTJ9WMf+Bi1PTyV
FkptWuITLpkYU4d54iuj1Ou1G4IOvsNJsEe1l0B6/q0qQdNgtnd4VWBHoVyrxvysBb5ArsmnJOyZV+i/oaVdyF7XVI2B765pTmcBEWRWpaosjH3S+4HJLLna5prva+NA
uDsaZBmMLNSOvjeWrjQM8E63+JORe46mAgbM0bdnmAUEVdKVch5YWxhoy8dyuHDtqXG1/QlYJTZ5JzllQwaI9k63+JORe46mAgbM0bdnmAXYakIzkXw3xDztKHbU+Aoc
omam5lLSAVTEeMZxoRrTFy0mycDcR7Lu0mrFjERaEAxYggDEwk5DWDzBxw7VtRF73eQyW3aGm7CasvYi55zkIc1hYJWTt3UUzZYpb//8FQ7T2qUD8KBDRQY1cIqQHL9D
6glR+5kww0XFKu0to/nGDijtv3dl28dzmm+cDUA/IaLPZrwyIw6FO6I2rvpxnoRViqzByd1YHr6IBCa17isjd3vGoJQ1WiUdvVpjSb+nj4stcTNsGKsq7XlETlqQBP/n
k4M1uiU8SJxoYU0pYtUpRi5wTy2wozi3+VuPFs63ZUf8mqYpKG/CFvK4v2+A6gUbq4AH5OudOyWNnCrJYzj5nxz7ocyWY6xBBQ2jUWsKP7R7/LeL/u4bmDsHy/iWApoF
zoYfLZYAuFy0nUG39oHmBuEHzoiDFtF0Xg01y6x5rvHGzIZAPMdrmxuTTgDjQZNnuY5z/UiHUqwsHvmOrlepRJBuaXujZnyxH7y3dTFWrYYdiU3Yfqtq64kV167j4YWF
rZY+XdSkH4lY6omSSWNTV5BuaXujZnyxH7y3dTFWrYZGOgj8sRYGBifMknTIGO9ABXHrW7Oo/J3hRT6snWR9NPvK6UoFI6JENGSIFUP2fJLgNywqiUGEQfI8nyI4ucnF
AieWUND8t41BAL1b1Ktw5fVmzVjn3i67DAmIcwasBWgvxSQcVNW/f0bJfEINWbh2vTRppGXLXiOS4d7nbmHg6N3kMlt2hpuwmrL2Iuec5CGwWip7t7P29mkuSC7gxY8k
PXHMYlw3k9AGhFIDJwtKOerWeb58Xut3tyAiW82Nct97xqCUNVolHb1aY0m/p4+LikWiSwEStdQMBFzF2lE1MquAB+TrnTsljZwqyWM4+Z8c+6HMlmOsQQUNo1FrCj+0
A9yTVhFmyiouSTkWdwXY3vWnvwvfNv02mp4sRUxZ24Wmxrdc9nBI97K7fCFNCdC6Vx1/f+kS1zVAd5GmTFwm2JJ1XxYpJ4CBzJILILhMHscGc9mm5iJ1om24EBZHu84J
h3tA+KOD+mavez+RqvOfa5DdT2rcUC5+gEQ/BhhH+/XRruXT0sePzV7TTEDVF9om6+mpT0YgYIjnJUBCj5cACt1fVzWxVY6oGOVpcEPXZTH51QxTKMrLBrXquCFeHN0s
5DE3yw8dnoNlWyoDotjqzfbeshtcbJO9GascshhESO8nkgUZPEKGvUGYacI2mVcxKx+1NNfqfV1FEw1Ul7QD5XJQo5MaQzs2o5PFuCZk/w8pQGl1wD9k+moe4aFzXIc1
i6qCfPbl59E4T9U0ypw7G+awyiwxiNkfP+79fkglyhmTgzW6JTxInGhhTSli1SlGLnBPLbCjOLf5W48WzrdlR4SBF92Ve18DamyniqYxO2DKiCbRJr2HgYyrX3ljAm2I
hc4jSwzDsq2W8fvr8FGgKl8/3zs0ko6wxwrBySYZspiHD5JyAnHHuD+f9ClzKIGEFkptWuITLpkYU4d54iuj1H0U3ppvrzO49isVRXPEHp8xYmf9TfvieZq4i1+4laBe
dALMNN7ShjAnyH1Pnkc1O5z1L2t3HIEPZNomGFGM4nMqQdNgtnd4VWBHoVyrxvysBb5ArsmnJOyZV+i/oaVdyE2gaPFuD+/VtrhBQgnp76aXkPFPtaUKFdsj1kx3zLx1
omam5lLSAVTEeMZxoRrTF0EoncHqtZSo8ytr3hQuwWTtWBYbDUTiBGknBSYu/JTYq3ZkKXXO2KKFUXqBJ0CXHjvtDHXdZZPhr/y9MewweBjPZrwyIw6FO6I2rvpxnoRV
iqzByd1YHr6IBCa17isjd3vGoJQ1WiUdvVpjSb+nj4uYRcGaJzxHYw+/jSMAXPz8Dw47LBKVbh0qT9gAJWP3+Rz7ocyWY6xBBQ2jUWsKP7RpdFed0TmriuqwqMxJGAm9
3tg36JZIjTN8D7VQ9R/Vso2F+Fy47p9sId0rF+e8ZPPkRp38mfMzD49jvGPw9yqaKkHTYLZ3eFVgR6Fcq8b8rFvv+mJR+f7LsT+qr0N0oEwpFzFsHn1YeK4ac44cds9V
gAdXtwqDtrkMcTULh34OFHiywh6Om/yrzO4ttzq6UeKtVZmxwUgP+z2KlEWdF6cuG+kiHRcaWrdZHDKG1hExGa2WPl3UpB+JWOqJkkljU1dKBJjz0YHOW7ryTJpxBaPY
IMYvlDvVq7PyYSF33tu4iZDqAv8LbHKLlrhNYS91Ol0jNMz2WdvGC1rtsWwsfqhCtCi53zskskiftcq1+bxinNdXALWgDvQVzL6zAfWYWZWzrQ6rdtIAjDaNcBxTnr2V
IFGa6Iewg4sel2IBGOtycFdzxTS1cBqmR8LtQuuJdEK2BLuVVekb0Xyl9Itst/a7PGnDdz7yZBhlZEZ79oomFdItQ2IfSpmWK8fMEo10RoeHhDRwQYb04w2mlavVwrFh
vxe0j5Y9NEHxBvb8pP6dPlGfKvss99kkAFlBAcwKnwZD8w3RxH1gqtnj8YxW9o6/V3PFNLVwGqZHwu1C64l0QrYEu5VV6RvRfKX0i2y39rvVKZY8BnW6/zceu3wdu/Uu
WqCk9ebz4VPo7nOqR2iEX61VmbHBSA/7PYqURZ0Xpy6pIwFQ9MHl/j1KoFBPm8uBi5IpdFCcD+FVTbzsNb9+2eWja0Jpd8UeIghUlIpSXBHbCrsFNtQlO8ygyYxdswGD
wnhpVTvwwoJr/ftGExDiE4euk0O5oTpSOFfwNZAei9QQ8uof69/eza0M+yJG/WVZBXHrW7Oo/J3hRT6snWR9NPEqhQUtWd47dYOx9wGI93GEO1LPhxGufbY1nrn+AM2x
7VgWGw1E4gRpJwUmLvyU2Eq49/KYrMzK0hhOkatEOrdXc8U0tXAapkfC7ULriXRC3etY48SK2ooG1Maanwdnrq7IJwfc0o2Lng6NZiBdODnbskS6rZvAxa5+jrBBT3uc
0HmRn8ralutiqQIzpdKiR721jSWOnkx+HKg0SkmdrkCBAgcgg5qKQ4g4aCbwgvbqiePltBa+MRI7/E/80opPeFmiWvqBLw/DJJb+4yfUZyhp9x/TVikdNR+F1KSEHESY
8SqFBS1Z3jt1g7H3AYj3cbVjndZ97K9Ai+1BkPzcyuiBkVhxHCywcQIJbtf2W4ygT4o+ycFjNLai+e5fFZWDz4euk0O5oTpSOFfwNZAei9S+3/HOMBCyzHRWLdfnEbTc
IeIg8YZdnTAxePyaHru/zSchNs4BkN0jWS/1+zhfKDxykdL38yBztMfrlRMRyQGkBHQeEgmFpU2V2oZrW8ortFdaHuRLua/3tZffJYtePQUXQZfR3pPQQxD9JE3WLcK6
nLZt7VhbFAJnvoCNP0w7EQf41bU2Mesjmz2xOrDp6UWclrpfpa5vo+0mlnRKikm1GUyhTz7s7mCobUZGZNbpgk+KPsnBYzS2ovnuXxWVg8+HrpNDuaE6UjhX8DWQHovU
vt/xzjAQssx0Vi3X5xG03GUvXig1hiXyhDj94sIVZvg1rkJgx2snt/UF/MNYFEAY9VhFLFQxd/SJbZjQr/xUvPg9B4LRSs33D6Zx4I6x4TDIZurXCP9+woMnU7RE7uCJ
R2xPEdIx7xRpEQD2z8jxgZJvvypUltaKxOKOZ7z2xvKiz/T6Tk7W4zOuo34YRfeKZzw8SoLjjdgHnAey4TmTOQUgWZRe/z4H7aIZBQyltdx59pzJjCaDpB2LDLHfU7H5
FXYR6m2Z6aZ0ZwD+pL++3PeH+oiUaKhlZHvCKpLPO8iLkil0UJwP4VVNvOw1v37ZH4Do5XbP5QRIHRZ/4BL+Oc75ZK4RrN0XbAjOBuhrJRQavhHwGe2ug9uTuSKoLOw2
9ae/C982/TaanixFTFnbhQ4E7Jvyj6b70G9yymiz4bZpWkNIkR52+B1lg04MPUyhZOPBketMLMQJFkuna2gtQfoiFHqHLUjtUhhvqeAmOo3+Zw5S0Yyrl0BAgXmSSmEH
+D0HgtFKzfcPpnHgjrHhMEgeo58QewtOkdJuLkdnIrJ/0KTxvCSFaxENyjQL8PhCsGQXNpsiZ5gm8jA43t4W1W3DGzAHATFJyRAQ8K0kHAIbfihAz7uVEbgyCGk4GuBc
xnEjtPpl3+NeCYMg1ynwNWeOmjt8ZM998NlGfHWRplnbskS6rZvAxa5+jrBBT3ucAVYnhivNzNQnNZF/62ZNg3dScausXeJ5hGascCe5vrTSTGeObs7fK9H/zE6InBQ5
1gmFhEo6zxk4sK0OCLzQ0ktg4j642iNd69D2hPjQPefdnFF/pAXdg6FdAIyt1HS9KkHTYLZ3eFVgR6Fcq8b8rFvv+mJR+f7LsT+qr0N0oEx39ESXTnGGSzLJD2Jvh67F
SfvjaG9uyRCBN4GOt7ThPsqIJtEmvYeBjKtfeWMCbYgfgOjlds/lBEgdFn/gEv450gqa7871niV3MIn5/MBvjLbng0xtNnld/dSELjm7j6lEjrhHO8pQ0unxpg8QWQMa
VovpwjX66oeTMs7V+XIbqFyPCbbkhFSGIDXrNVtHiZN3NhFJimsRasEAGHoikDVHWeYpyahGuqOZ5ZnW61KVN8HGuSRZBeQ1QlxYdvj3E5idJmLLWuxUy50ApYJNJjWp
DT2KOrsT9gjx9wo9umnRP5JvvypUltaKxOKOZ7z2xvKTeoK/U1PfG0RG9guV4H+PSEE/RIUPM/uKy+F7A5BNIbmmsO0xWGId8kQtyhwvlp3COv2nPumNChLTfqz7pfxg
LMX0D9Mp4Wb2ZGI3yRiJ3p8cYdZelJOjvPRmgkiwPTRWBg2q2AiZrAIew0p8jy1p3DJUyJbFpI8kNy1xDzzcT9uyRLqtm8DFrn6OsEFPe5z17ET+DYV03lMnauL4fHAO
YswXAGLSPoa1xmiwYefboQ09ijq7E/YI8fcKPbpp0T+Sb78qVJbWisTijme89sbyk3qCv1NT3xtERvYLleB/j6qZqlinSfcSiJ+KmLr8CWxjhG8JtiZjrwROw/MW4NQv
uOMB16oyxClll7YmYnuL1kVWYGeElHmQyIv6Jf/sZMGV6G30YF1NLY8L8JbTtK5SKkHTYLZ3eFVgR6Fcq8b8rFvv+mJR+f7LsT+qr0N0oEwCRuNiT6px8o77V6Ex109Z
5Deb+BY5FsKqD2oOSLwiG9JMZ45uzt8r0f/MToicFDnWCYWESjrPGTiwrQ4IvNDS8mOg4CWLLsI4RMaIXEGyMMmRPHfzMmq4uJ5FmJSUg2G9yeGw3O1Gy+fHoQQxwBTC
5j4J8UJVVqyAilSQiPlR4x987aLTnUqU5WBDSxbwAsdIHqOfEHsLTpHSbi5HZyKyZWjMxhazqdRPPJa73fmj+VqgpPXm8+FT6O5zqkdohF/hB4i7RFNp7oT7X0hIxZQL
cimFcnn0/m00dAxHyTVa4e3W5iufZM6wN+8aIXbsxUog4bhbVoVNR8l5+tmh9qcWSgSY89GBzlu68kyacQWj2PUBvRbscYGJTTBpls88kX3tElv/2Q6e9RLtFMBalWHU
uTokCP30q+mI8WpvbNwc4AYCTeHvWsY7j3HqNqNoCspFVmBnhJR5kMiL+iX/7GTBFXYR6m2Z6aZ0ZwD+pL++3DXRcL8e15Zs2WhMrBcQsKtJcGXfE6wIoe5d40MdW6Ra
hhhVdkMfQzUMgopFUjH8SnjqFcViLTojVUaaO51H3OZlYNgUgDVcEjiOk+iVgCyiHQ5w1eFb0JYTrKrbUeNY5oeuk0O5oTpSOFfwNZAei9QMV7GKYfAi6dtC+Zgv/uO4
8aueeDpm6fRHb1mn2YrYvzWuQmDHaye39QX8w1gUQBj1WEUsVDF39IltmNCv/FS8LMX0D9Mp4Wb2ZGI3yRiJ3m3nEkl1ZsgvDyf5WfWldeCQ3U9q3FAufoBEPwYYR/v1
1FIXRCphps/WwxNPouZdD9cvhkaCq4B0ohHxWupwAz1qdaVJY3ejJ6yC+HCzYXYI2cG047HjYtqQmuboNspyZSQfIuaNjTPke/SdYEjXTxtAVflo6aiYwjAHv7TsxsK3
bSIGEXSwPhnT3DgKa9FG1eGdkjlIuQvKjIu+stmKKZ15CjPuutR48as7YARutKNFLrsIHtNO4lu7EivG7v8spnKbOMRcCvOPfekKKFd8kK0SPdVWOOBiBObQxBzoIo1c
fZild8l8Rar7/p1EWrBHxEvVV7b0zi2pcb6wLohqRbSsKlkRS+PAw8OV9jhA20vo5MTHwCPNcns/aMRXjDbE3v5nB/hLOoJ/zPdgTOGFX9Gl+hFDaQi6whSctnD6VO1w
t4tonZ/uPsgF1gg/bcH8q8apZCQExvPmf8enBuf2aS0mz1UfwqE6SQ60Vv7qCLXOfHqotDeMknfVw46sdxMXwSg5RVvHHMh21YviZA1YquAzjl/3KNjeNMExa+jpN1e9
GzosaODw1bolQv/E7SWbpbeLaJ2f7j7IBdYIP23B/KubPaaHFZlcNowvMdFltcdFNtXnXeVzf94QRinks/40Ec91J5lFGk/mr/CWsyccKmpNwyXsaEasSuMuLIAh1w9A
ZbDO/js5xZrSK8JEzMQCuwbGEFSAxRjkkZG/BQmmxtZtIgYRdLA+GdPcOApr0UbV4Z2SOUi5C8qMi76y2YopnVvlB2jPPT30xkvduXyZqXSL4NuL+5+yyNvFPwb/TQKK
KolYqjzXPXDaBXqtcyVsW577b627mK+HMiFYzz0LpL26lzXiAK88LJHwXSazsT+NdKq0UrKGIWMmGOapl9lvjEBV+WjpqJjCMAe/tOzGwrc7ovk4t5Ol47NGJvsKX4Yv
sLugnDhjUR3ulT5OO27Q9Ez2kExSniwT0lI8sasg4QvKiCbRJr2HgYyrX3ljAm2IEt5KvyLJ2M92v/NEKJlk+3c2EUmKaxFqwQAYeiKQNUdSaM3YW+iOYEhTngayst1r
wbyedZlwNEf692em19x1xcqIJtEmvYeBjKtfeWMCbYhz+zdJoLhTmOCtgEjRTAYGC6A5qpX4zaD9YzP3omMO0ka60lyyCjM4zjOwd00CEQN8AbGimwFwvtzhog+aXy4a
sY0fvbSNx0+MJqfNjmpwSdu6+LDvqdi+9PkQxQs4MvIBiXo8hhvh3EmXU6N8/btKkVxrQOJrOZsrNtfakjOOGecNmYSRq82IfYhMCvE5fXosgXLyjncDCJdbSJ6UpwT8
gGKA/EzuNW5fsOqWypwEs3TBiDZG9if88AY0oQjnFcYUkNtLIYtdFhC7CGgWuf3CKkHTYLZ3eFVgR6Fcq8b8rKw2+H+D/hSMdX6vlX7WClUBFrVPPqZPd4+4JZzI4Fv5
dMGINkb2J/zwBjShCOcVxuF5ew+v8pOut+69vGH7iyGSdV8WKSeAgcySCyC4TB7HeUziShtIZ9jQ1WNWaV2RdGoFHXu1ZCmG3bhV3wbEcCFMk7aOs58AkAS7w4D7A0lz
RuKJl4yWeyXU5zcOzNMYHwP9bEmm7ptGufiEOwjFk0r3fFiltSDf74ExyPZuc8BOOiPMB4BwZuzQdZVhDLLIFcakdCWPm8GRN5J2SM4b+JKf+GkfYiIalMywY3yWE+3v
O53DZpJaBNjYpM9WmnHJJQ8kxWRPpKAatSVRsRjAsz86I8wHgHBm7NB1lWEMssgVlKPloq5LGBaG+UU3SRTQwLv8P6pmnBvuHpQN5LO0jdC8D5BxaT86gUjhxRmy/L7T
H1eBs6KoH1yFUljSVIl01sqG60/noq2x6qwFAg8xJXNu1NyM5fwyusOGAHmWwwq8zwL9oEM5mybydtbqSNOBiE728kUeZ7sin9oWLIVFvlNL19nAGIQCD8bB3Gd0DFv0
DPGJ4LlztRgXXDfIuFQsPYvKvqUAxMn1Yx/4GLU9PJVUKnn93PYqTBxtIQwia/aF2/kCIcUfW+/KLSRTCF06Y7DPrCzgt8ho6MTxoAaPvYnj/FBmgeSPyUOFuJvPDLWm
N66FNCoreQ7Y3+8bVYv0SJJ1XxYpJ4CBzJILILhMHsfj/FBmgeSPyUOFuJvPDLWmYL3vMpjZA/eO2aDmjv68BXYVFXW8Ph0+MM7ygckdEfICoVYdikYZemG72u9hXwCr
BxgFsQG8uRW5zXmQOf61TsqIJtEmvYeBjKtfeWMCbYiyqwpkE45yFXuZv+8M/oe5TwwO6Lm/fG1Y74BvtPpzDwKhVh2KRhl6Ybva72FfAKsH0QM+dk9wYutxNz1cWQYM
z+0K0iYUMQzQULqZMhffgXSKBcpHnZK1lS1b/PV9NAhKlCNmEZGVUT8wQ3TXTdnvUQ3RcVVLuo8f8A/DJ0FOsY4Qwrb4q8WTg2Jge60/0gs/GTU6I7W/A6NjnD3jSmcH
0kxnjm7O3yvR/8xOiJwUOY4Qwrb4q8WTg2Jge60/0gupeCERDt5oi3A0ohoUGqLAUaLwr5BdD5vS5yulP3+e0w00RX1Czr4bLJtienk3Hcdh4YAPvw4jNAzwO9MVn5FF
JQIN6+P0OMns8Doq3JiZIBqUom8LPbntWSHX+jZ8NcrCeGlVO/DCgmv9+0YTEOITxQXWjVoY8rMqF0yahEr4P4AHV7cKg7a5DHE1C4d+DhQShKruXmOJqEJC4GCzlmIy
aq6wrekiVqzz5hDbugBn2gugOaqV+M2g/WMz96JjDtLPlWvvQaLR7ZKedRBT4OyvrHDMgBhvE1o4MEPqMaxIwHMl/QcigG+SxjraxpZtiKcTr7fBIMYTkjBP05A0/fdG
u9wut8dIIX6I9l1QxpEatEqUI2YRkZVRPzBDdNdN2e9RDdFxVUu6jx/wD8MnQU6x/s2lNV/hdKU7hL8BqtLZfa4WVpCiBDWk3zRHo1U5q6YYjfA1VIJo4cY95FP9oxnu
z5Vr70Gi0e2SnnUQU+Dsr6xwzIAYbxNaODBD6jGsSMBe6EkKgv6tlb99kI4RmTrIq+sAwRY84H0iuscNnQ/RsbvcLrfHSCF+iPZdUMaRGrTGcSO0+mXf414JgyDXKfA1
QNyz0ic7B9l/jnbp5O/gyVssvp1rTTekVeHxaqbXTIFlYNgUgDVcEjiOk+iVgCyiT4o+ycFjNLai+e5fFZWDz8UF1o1aGPKzKhdMmoRK+D9gve8ymNkD947ZoOaO/rwF
dhUVdbw+HT4wzvKByR0R8tWnNbKGYFVshvdLH7ovnGospSLROrGetzsRP1bFobXaR2xPEdIx7xRpEQD2z8jxgQTGIDLjVMJsv7urJaPnSB8BFrVPPqZPd4+4JZzI4Fv5
gUvN5SjjrElx1qGpcAq57gNCUql16CO1fFB/dmWiAxp+q2MKRnK+BNlMXYdJl7zGH8pEsnRSHrYQTi/92R7xmjiHe4O1iAvHhN3WGhD0oUndDxOLItr8uVdUPS31nd2R
nmn2ungrLgKNDA3+nL/zM3y3H4EPCCVughaBoTnJXSfjSrvr0a/YmP9XPo5lFoAuVuOw95SQO/1Q7fKPYfQLnFTfP8zuuwnXLmbDJX6mfuZhsWwLXHAoNbyYilpKhZNl
knVfFikngIHMkgsguEwex8B9QFnD+bWrMFvtMZqlYL5hFvMjZAIYRjUP6qbaWioJLVzyL0eTV5i8SMk7EIMRRNHlKFEiX3hS8GwLUzkUmcnLi5w5Ul0/WqA5tMBlxgFr
z63Zoh84o477Hm43Km/ZSIAVFwoUFuI5PVf+NIlC2I2orqXdKFuVZY0h1osc8y5S6zzsXpRNIxI6RaHrh0RcVY3r3bzM7n2Lz04uEcMWtTJhUqSvC6EjN+JM1BloexxE
/39jK1a28UYbNFEZFWPn80THtIO7IXRLkgBzXAaIVwlNCCm6LWRKQPT1MyUfei2DQ+GzYUPcEjn/YlLkoeK3s7r/d6zTt+cL7zyOVXqI7NBhUqSvC6EjN+JM1BloexxE
dwIft1vyZ+O+nrvStz9g++hcrbLYjACUujisbOLLPEiTUZmc6FjBEvPzR9vujdoaBHj1g91rCwqO5hTfLniW4B0OcNXhW9CWE6yq21HjWOaTUZmc6FjBEvPzR9vujdoa
lYw/RDcQlIngyXzd3C3B1yhUcgoxtL5qmxVnrMJ7+6Z8QRVMIQ8kC3djBy/HzmKTs87bwxNr91TwlIL3efE0+JJ1XxYpJ4CBzJILILhMHsfa+UkFoverjWWKkUZKcSsn
2aj5zAlvLkIcbTtEImNHnLSi42CibOM+/jEPGNo3WyO7EcAKVayMOaPsik3jKbDdJNCAZ56RmEDFM3SpohEZpwjj8IH0rH8pDaqOV727uhquouzwdWtjCt9owoXxE5Q1
APJ1vJZcTF1YQEMxWNiL+fjbgiUqlrA5YtkrHcOd8EhhDbrYV1Ft1mEAQ9QJlHxxUaW4fX2pBEJnZuYqxpkCaewGAYFmU79MPPKZ/tz4nGXrsK1wupmEpoCynz/bdPSg
MC2CL4FJQAlZEkxpfmhVMe1YFhsNROIEaScFJi78lNjR5ShRIl94UvBsC1M5FJnJJPh677B2YLRwYWFiUQpraArjUhoIMMVclD6PUVEARyvR5ShRIl94UvBsC1M5FJnJ
JPh677B2YLRwYWFiUQpraL21jSWOnkx+HKg0SkmdrkBVTFcJNWYysVpHtG7kevqGJPh677B2YLRwYWFiUQpraIN/qRvhWwjvKE0755rKsOvwTHCwzEObuPwhSv1lPYL/
xr8CK3RD+7d7egvmMSIYGiO4BkcxQCmgii+ZVhwjczbrsK1wupmEpoCynz/bdPSggZFnmeSUE5RbnedElXMLLaoO8NN6LFd6t/5dovnm6IjKKNmHwubB+IqJtf9aQLJk
sVeZXS2dbIYw2f976oZSmHc2EUmKaxFqwQAYeiKQNUfKKNmHwubB+IqJtf9aQLJk2Vgcg1FIKrSJTHewx6Tcwz1kguzPMN9cBhhGj13e9piyI55EoEIEokDNjDUTCb95
2QergHaszq/6gS+1RVOZ/6dNG2tI7fwxIiuSthHusS8xLFNhjd3n4e2W74alQGlSqK6l3ShblWWNIdaLHPMuUsvCUc90x1uyyIqzT3Pxc1atlj5d1KQfiVjqiZJJY1NX
czOnC534/bgvwa0RypMZvcdqVb00tQYA/JMP/5wI0Zmtlj5d1KQfiVjqiZJJY1NXczOnC534/bgvwa0RypMZvd0Ywdm4LNUDmS/KYJAyybP4olUzT5ombdI1SbsmTTeS
voNpBvkHMm+pybjOlltiOJtdX/bTGsFaVlQfoDpC3WcoVHIKMbS+apsVZ6zCe/umfEEVTCEPJAt3Ywcvx85ik0mh5Gd6Hn1Tvv0a4RXA3lFEx7SDuyF0S5IAc1wGiFcJ
TQgpui1kSkD09TMlH3otg3le/4p26IM9Jogie+SdAVjcD8/GBBhaBgkLK12fVWpRYVKkrwuhIzfiTNQZaHscRJZUahi//w3LNUy8rHd9FZbkxMfAI81yez9oxFeMNsTe
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mODXevbED+b9FmV7bUbifGoKkHTYLZ3eFVgR6Fcq8b8rAfFtt6jBmZr/DhVrKZCJx1nckI1i/bOzDo7hjcWHXWn
OZIOaATV5WaZ0+/AUfSa+pS5hx1E+tr0pjHaWfBf6rnsVU3OE2J7ycTS0x0spYZs0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mOumEc6sdtfL8qTdJIlcN31
KxmX1OGAzUoDy2epYk1OYjEsU2GN3efh7ZbvhqVAaVL/quZ2O1gb9ksqyxwSuwFISNZodRTQofIbQ4VJyf6YGbyAJlbaCENd2xijg8aRizpp3lo0a1J0hEzy2LVT83uo
3Y+e4YTMDjyZicr+JJtWH4dZlUU3ULhl2yql3ESG8Rz/w4vxX/mfRPtiUY9y2S8aON7OPUdOLajaY7d0vFdbz9gbzrfaFm71ShrXlUko3L+EQhAYrTJaeyyfJDIreORK
tpzsxfRgVAH0LvQCU/Sx12j9cy7XxalrE4vLfskOs3rOMywmofQzuM5YrRxCFA22tYFtn1istTRgz5rEHLuDwbMisVzkHDO/pw0MifpxxA3WQN5NBJ63YRSJ8xjWyfzc
n6idFNTjcyGdFocxjFlNsiTi6Wul/Hh+DEXd3GiTTT40Txg9v4IN/xsDwjDwe9QusiOeRKBCBKJAzYw1Ewm/eTRi6/Q7+mjbCiqWtUGmNqwnpct/UjXD7BYTEByjkLBm
owOdxnyGU+bJm5Xykh1LJX6rYwpGcr4E2Uxdh0mXvMZo2MBLOkM3JW1YJuk/IZ/CNGLr9Dv6aNsKKpa1QaY2rCely39SNcPsFhMQHKOQsGa33GsaiXtXsZ3EqlwkGBZa
72p5AS3MDP4vRGP69joIc0gYkj1yTntkFNGBfPjz/LV9RShOX4pAd5/GmofNusGv8WYCQOe3HM2U7TOn57FjPAIGrUVJnUR1t158n7nXQbtMk7aOs58AkAS7w4D7A0lz
SBiSPXJOe2QU0YF8+PP8tX1FKE5fikB3n8aah826wa/xZgJA57cczZTtM6fnsWM8fFGh8NBx5umhptrb37Kuy5s8e8iOIgREIkjUYfkE/nuWPtBTUaG5LS29LLwcVRV/
/cORsL++nfNhMApynjsK41wyIZwcuUxMIfE7Xw7+GaYLW2X80eFSwqdlbBCXyCEGrZY+XdSkH4lY6omSSWNTVwcz/AzImCCIvXvC41biajt1wLoUYjnAAEjwaCBgCZ6K
AQVYFhZzpR7XPEeXoFshVcHwQRHloHr0ZuWr9vnWpmlRovCvkF0Pm9LnK6U/f57TBzP8DMiYIIi9e8LjVuJqO3XAuhRiOcAASPBoIGAJnooBBVgWFnOlHtc8R5egWyFV
eeZQv7xEuJVV4PgeIXMOFuCsCD3UlWynLeS4fDBjEsb/quZ2O1gb9ksqyxwSuwFISNZodRTQofIbQ4VJyf6YGept5fYFgXGhC/j93uCfMHGMhoU3uKDXFb6Fj7vx5sWt
UDq5J8lZxFgC9xYjbv2iAIdZlUU3ULhl2yql3ESG8Rz/w4vxX/mfRPtiUY9y2S8aTC3RL8uUMQl2nzsYuvtERO92pP+koWQ5dxWSUcIA82SWPtBTUaG5LS29LLwcVRV/
/cORsL++nfNhMApynjsK41wyIZwcuUxMIfE7Xw7+GaYNtBuY7tl5LrZoPAfEtJme4dcpIwTJlD/fNvowtATWpQcz/AzImCCIvXvC41biajt1wLoUYjnAAEjwaCBgCZ6K
AQVYFhZzpR7XPEeXoFshVbXGrZljn+hZzjMcgXm+d52Qf5HmJoBE6WxV8oGBLTtqq6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCF8hCHDjVOli38TUVLit3RG
Xqe+r4/CO/CI2/Y3d/XR6DEsU2GN3efh7ZbvhqVAaVL/quZ2O1gb9ksqyxwSuwFISNZodRTQofIbQ4VJyf6YGept5fYFgXGhC/j93uCfMHHp6MF+MoRs/l4UtyfmKb3V
T3xlvNQSevanAtACsZiuqbac7MX0YFQB9C70AlP0sddo/XMu18WpaxOLy37JDrN6g/rUGbM7MuzAcC9OGCPGpv37JpZeAcVIGozBl5NTvjiuouzwdWtjCt9owoXxE5Q1
NGLr9Dv6aNsKKpa1QaY2rCely39SNcPsFhMQHKOQsGaKIEh+RkMVD+zG+Vp12EzXD3n325gmAMc3/imIJPP3av8V+cqXC4OEaSDMT0wEx2xnckI1i/bOzDo7hjcWHXWn
OZIOaATV5WaZ0+/AUfSa+uF7a3IjpcSsS7xYtBfj+or8L99vaqKV7jG9Lm8ARMTP4vxlw9YuKkvFwCnfglX19g5pQuUrhjkblzQeOns6JP6eMbn4yOgdIHNpsoDnqgNH
rgOoFtTixhm3zEBZG2GN4NwPz8YEGFoGCQsrXZ9ValE9MI5bQvq0DRFT9Sp/3zYuaY3SecHz2Z+yApnqIuEE+BClp6dUK/9xWmNfz/MpCWiuCiBkDg4SQZLfoJnJX2E9
gBUXChQW4jk9V/40iULYjf+q5nY7WBv2SyrLHBK7AUhI1mh1FNCh8htDhUnJ/pgZsuGgY4ulq2aX2YKDLM1hI7Tox8EJU/aayvfFx5bXxCbkxMfAI81yez9oxFeMNsTe
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mNSTRej+I45HK0oqC+8rtFuvIE6JIR3wvmDGvu6AO7ulY3r3bzM7n2Lz04uEcMWtTI9MI5bQvq0DRFT9Sp/3zYu
aY3SecHz2Z+yApnqIuEE+GbpryntX7HwLHo9PhKV0X69w5Wj2C2S2Ta8yO91umlrcFZfXSWvI+nGKVpcfce8gj0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4
ZumvKe1fsfAsej0+EpXRfv3KXbzzWgjRzrCGczMJsyC6+9x0TU1U+1qDZgR5SMhe/6rmdjtYG/ZLKsscErsBSEjWaHUU0KHyG0OFScn+mBmy4aBji6WrZpfZgoMszWEj
nzMado6RaLHuOznH/TWzMdMREg7XYI5gppsZMW1kELE9MI5bQvq0DRFT9Sp/3zYuaY3SecHz2Z+yApnqIuEE+GbpryntX7HwLHo9PhKV0X7N3c+AsJ5nCPh3iArsgnMO
na3GG+kmLQjH8phP6rfb4NIGiqxNdkF8pLgKpY2b/XsGhtgRD42HToRY059LAeJjUk0Xo/iOORytKKgvvK7RbuRvss3MI6IX0eACanheVM9t2hFLlc8LQ/Ink0BJ0rea
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mNSTRej+I45HK0oqC+8rtFun/OJhfwq3pKHya662RAmnc0sErjYpIovT97sYzYP+aU9MI5bQvq0DRFT9Sp/3zYu
aY3SecHz2Z+yApnqIuEE+GbpryntX7HwLHo9PhKV0X6O9Gz/Wh5L2B8j8/y11fb3uv93rNO35wvvPI5Veojs0D0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4
ZumvKe1fsfAsej0+EpXRfkvuVb6F/OACmJzyWXzoWDjmjYZGTPpx5fHkDH12aeTGq6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCFqyK88yGeJYhmhnXyR+ITR
H/snGXyui588P5S5Ff9NlRuvFwZ7uF76p65+MYtmN4g9MI5bQvq0DRFT9Sp/3zYuaY3SecHz2Z+yApnqIuEE+GbpryntX7HwLHo9PhKV0X7SsvGUUDSHAePIh3o7r5LI
3A/PxgQYWgYJCytdn1VqUT0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4ZumvKe1fsfAsej0+EpXRfmABSPr2srLCLVgIC6ejzZ7KiCbRJr2HgYyrX3ljAm2I
q6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCFqyK88yGeJYhmhnXyR+ITR3WGp1YV48LbSwTfm6RauUyfZcsbr8AS0IXcujMUDRifi/GXD1i4qS8XAKd+CVfX2
DmlC5SuGORuXNB46ezok/nVzWclE087CW6WrMnOpGN5sly1X1LKwUvNsn+h0ez+HqUQlk8qqei7ue7/eaZic1rIjnkSgQgSiQM2MNRMJv3k0Yuv0O/po2woqlrVBpjas
J6XLf1I1w+wWExAco5CwZqikO8XQ8Bb78lzeeDnZQ8svMRcRU0wFs2T7MxA7CRed/ozHgkCqtaWGn4lSW4utgJGlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKU
OphwATLtaA5C0EoIoK1V9A20G5ju2Xkutmg8B8S0mZ7h1ykjBMmUP982+jC0BNalBzP8DMiYIIi9e8LjVuJqO3XAuhRiOcAASPBoIGAJnooBBVgWFnOlHtc8R5egWyFV
IqeLZk7r7eua92aXU5JOxmGBI+kEN5wAnqfWiQJ/QXmzIrFc5Bwzv6cNDIn6ccQN1kDeTQSet2EUifMY1sn83J+onRTU43MhnRaHMYxZTbJKi+nm/VD8hzx4aNJVIfHk
wxGBydeLff/vEf2iiACq4XBWX10lryPpxilaXH3HvII9MI5bQvq0DRFT9Sp/3zYuaY3SecHz2Z+yApnqIuEE+GbpryntX7HwLHo9PhKV0X5ZQv+Yh/5IcGX0vCUhMYge
Opeok1I1+qBzUkkSmfKCLP8V+cqXC4OEaSDMT0wEx2xnckI1i/bOzDo7hjcWHXWnOZIOaATV5WaZ0+/AUfSa+rtuz42U1AXkK8qVYyP7lh02fc7IB6c2eFfJ5B8M5eAw
/ozHgkCqtaWGn4lSW4utgJGlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKUOphwATLtaA5C0EoIoK1V9N7//AtJdwzYO9hTxOAMkToiGP8sbF0njmT7/2yI8rkq
4cxe+W8T1i50iFuqTkMY0P9aPE9sH7MI42fPI4d1a3m/bUOMp9282Mxd3WcLOGjnVIJ3CHSqo2a/BkQFiXgtl5SwoyToGZxVwvAs1PhB/l5hDbrYV1Ft1mEAQ9QJlHxx
NGLr9Dv6aNsKKpa1QaY2rCely39SNcPsFhMQHKOQsGaopDvF0PAW+/Jc3ng52UPLvvTXx32PFCa5IlixsDvrKuTEx8AjzXJ7P2jEV4w2xN7SBoqsTXZBfKS4CqWNm/17
BobYEQ+Nh06EWNOfSwHiY1JNF6P4jjkcrSioL7yu0W4LsQrSBZJZ1KOa1r2riUOOkN1PatxQLn6ARD8GGEf79XD+hC8NPCn7/nGyetCc8aT9w5Gwv76d82EwCnKeOwrj
XDIhnBy5TEwh8TtfDv4ZpiO89ehnae4HfBcjsDToaODtyUsOJD3CS85a7SzIsCE7y+/KBcRvy6e+qn/l5K8lCodZlUU3ULhl2yql3ESG8Rz/w4vxX/mfRPtiUY9y2S8a
w04ZNB0m27sv0riZEJG8aYe94sgwcr2yPz8JOfh0yhWN6928zO59i89OLhHDFrUyPTCOW0L6tA0RU/Uqf982LmmN0nnB89mfsgKZ6iLhBPhm6a8p7V+x8Cx6PT4SldF+
cCiEixG+5iou7yQmj6w7vihUcgoxtL5qmxVnrMJ7+6bhzF75bxPWLnSIW6pOQxjQ/1o8T2wfswjjZ88jh3Vreb9tQ4yn3bzYzF3dZws4aOfe2m5e9Fboi3XU9lsHWDYW
sM+sLOC3yGjoxPGgBo+9iZY+0FNRobktLb0svBxVFX/9w5Gwv76d82EwCnKeOwrjXDIhnBy5TEwh8TtfDv4ZpmwTJAS3Wqw8zXCbweLr7x3YG8632hZu9Uoa15VJKNy/
hEIQGK0yWnssnyQyK3jkSrac7MX0YFQB9C70AlP0sddo/XMu18WpaxOLy37JDrN6QLfcNwWVyqlTPFJKx6pcOeyPrpgHGugW6zYeLLlutvudrcYb6SYtCMfymE/qt9vg
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mNSTRej+I45HK0oqC+8rtFu+1l0qxjGpPTqDUKuALHN1yt4yzJRwMwbtPp+vPYF5BHi/GXD1i4qS8XAKd+CVfX2
DmlC5SuGORuXNB46ezok/nVzWclE087CW6WrMnOpGN41JyqBcAns7QhIyk8PhxOGC6A5qpX4zaD9YzP3omMO0kgYkj1yTntkFNGBfPjz/LV9RShOX4pAd5/GmofNusGv
8WYCQOe3HM2U7TOn57FjPK35tuZ2cDJhs/rmDp0NW3ujZ+4MzfLK/DbXPiSYSM1g7DFhx+bklAnVUt7ltfN6fbac7MX0YFQB9C70AlP0sddo/XMu18WpaxOLy37JDrN6
QLfcNwWVyqlTPFJKx6pcOaUi1wQJOv0cUcfmb2urQBPmjYZGTPpx5fHkDH12aeTGq6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCFqyK88yGeJYhmhnXyR+ITR
jwtl7CsCnSGCnKP10VOXJoEhFAYoSae30I2gFsc9QvLhzF75bxPWLnSIW6pOQxjQ/1o8T2wfswjjZ88jh3Vreb9tQ4yn3bzYzF3dZws4aOfIRvPy8ED0V5jyYakDha/5
YeGAD78OIzQM8DvTFZ+RRQ29QjKh5tOiuQYB0wXkQkN9RShOX4pAd5/GmofNusGv8WYCQOe3HM2U7TOn57FjPK35tuZ2cDJhs/rmDp0NW3uhbpR1e3qhZeRTqoR0l+2l
mgYJrmRJAEoOTs30HnIF5pGlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKUOphwATLtaA5C0EoIoK1V9G03wx7+M1C6qYev7rvmATsn2XLG6/AEtCF3LozFA0Yn
4vxlw9YuKkvFwCnfglX19g5pQuUrhjkblzQeOns6JP51c1nJRNPOwlulqzJzqRjeIrSdQm+FrShaVenAAMyR3uPg2L1PQFCgMLFN4MZv1wHViQAJiX9c+A8e1PgmbvXA
kaUI6BdDB4cBakAqvDTW0srOfndS1iyFM5PAOFIyQpQ6mHABMu1oDkLQSgigrVX0LCrisFimv/69/+dSe1m/TiFI9tBXcYOSjEk5I3rXDacHM/wMyJggiL17wuNW4mo7
dcC6FGI5wABI8GggYAmeigEFWBYWc6Ue1zxHl6BbIVVySQ8wX66oevQJVCSgePlpBOYYhtua952DlVIopRjMWA2qE/AP1FXLbo1NuuPl8EWrpY9OqzrTG3VR9UcCk3LY
nreOuqgKTuhm8gA8sOhYIWrIrzzIZ4liGaGdfJH4hNGNGa9fO6d6G0QgnRcpiWxKYYEj6QQ3nACep9aJAn9BebMisVzkHDO/pw0MifpxxA3WQN5NBJ63YRSJ8xjWyfzc
n6idFNTjcyGdFocxjFlNsmZovmyHAqJS/dqDd4iuSMsI6mVnIaic7c40PQK5py8XnlzQW3r11+RaB+HzLkTUDOHMXvlvE9YudIhbqk5DGND/WjxPbB+zCONnzyOHdWt5
v21DjKfdvNjMXd1nCzho5yjqDIb+0MnHhCtZVW9pDluoNElbGaFvTPoyyBDUrL7lB/ypdMCixTM+lioGCXdQxNIGiqxNdkF8pLgKpY2b/XsGhtgRD42HToRY059LAeJj
Uk0Xo/iOORytKKgvvK7RbjIW/3NuwwNsSTGWpKVMYID9+yaWXgHFSBqMwZeTU744rqLs8HVrYwrfaMKF8ROUNTRi6/Q7+mjbCiqWtUGmNqwnpct/UjXD7BYTEByjkLBm
uqjgxVrQj29G58UtqHx7rBGL2VeZ0RNKkSrZlfI7bj0iGP8sbF0njmT7/2yI8rkq4cxe+W8T1i50iFuqTkMY0P9aPE9sH7MI42fPI4d1a3m/bUOMp9282Mxd3WcLOGjn
KOoMhv7QyceEK1lVb2kOW/oVm3mIB9QSYRtXFVEZ6Orm2yqwPjlNDdnx18xVZeeWkaUI6BdDB4cBakAqvDTW0srOfndS1iyFM5PAOFIyQpQ6mHABMu1oDkLQSgigrVX0
j8UaVMW5g7Kpi84pie/+Rjlrf2hXCVN1zEJbu2INdUwHxbbeowZma/w4VaymQicdZ3JCNYv2zsw6O4Y3Fh11pzmSDmgE1eVmmdPvwFH0mvqjfsWuKq5lr+IihlDWJbcy
Dgx9KUYLi+SXCYizfDXaa97YN+iWSI0zfA+1UPUf1bKveyi0N13qZ4pHIXwmOETsel5Y0Fv8O2ddyK8G3ChpZ0qxoqsLOMoQSNvg8VtjYmVp9x/TVikdNR+F1KSEHESY
Db1CMqHm06K5BgHTBeRCQ31FKE5fikB3n8aah826wa/D7bkaZSjg31gI9RJjLKxUZu57g17tbF8FcoohXgWVjrHuBmMjfXJGAqghOrGAz2P/quZ2O1gb9ksqyxwSuwFI
W7z9J3VFbg6BYeC4mcQjys4zLCah9DO4zlitHEIUDbaDf6kb4VsI7yhNO+eayrDr8ExwsMxDm7j8IUr9ZT2C/4dZlUU3ULhl2yql3ESG8Ry6N+d/wtCY92VICekCyBqn
lXpWb0YR1W5aCpYrA5R2NzPEOW9l12ScTCtyYVqrwQoNvUIyoebTorkGAdMF5EJDfUUoTl+KQHefxpqHzbrBr8PtuRplKODfWAj1EmMsrFQKZ46XNL+6lZHxiLR+32/d
UaLwr5BdD5vS5yulP3+e0wcz/AzImCCIvXvC41biajt1wLoUYjnAAEjwaCBgCZ6K4LM3LXag3oR+bD/1mvj2/R8e65sD5Gu7Y0bwhuyPVA1VTFcJNWYysVpHtG7kevqG
tpzsxfRgVAH0LvQCU/Sx11jPGARlgPg/3/jJcVUEG05a1cotR/7h5K6DISbHnbWFEZZspM1sVJqBnQ29OeFIGu4HofXgcH2cyPJna9UBQ5JnckI1i/bOzDo7hjcWHXWn
2YPBqGtfW5kk9tUQ9aDUVJy9u00+1gdDiz3Jj3wgbpDKiCbRJr2HgYyrX3ljAm2Ir3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWcdglqrDLQbqsf/8CsoUl4Z
5b7MF6tTq5i7Bg3yznsPOZoGCa5kSQBKDk7N9B5yBeaRpQjoF0MHhwFqQCq8NNbSccbPsU7g7sbfjv237YicWMNOGTQdJtu7L9K4mRCRvGkK41IaCDDFXJQ+j1FRAEcr
0eUoUSJfeFLwbAtTORSZybac7MX0YFQB9C70AlP0sddYzxgEZYD4P9/4yXFVBBtOSovp5v1Q/Ic8eGjSVSHx5OvtgYcisHDv1lVcwx9z2M/AwwEDDR24tENsD2/Ij4Q5
h1mVRTdQuGXbKqXcRIbxHLo353/C0Jj3ZUgJ6QLIGqd81oTUjMIDbjD3blvkP/iyTxWQTlI1C8BjUyKHzBoZ4h7w5HH6GboNGvHLqFXrEeo0Yuv0O/po2woqlrVBpjas
/uHALr0mP1efAQxMWRjDbJIDyVgPwzRAK07OJRXuUL0qQdNgtnd4VWBHoVyrxvysB8W23qMGZmv8OFWspkInHWdyQjWL9s7MOjuGNxYddafZg8Goa19bmST21RD1oNRU
hOYdZ6sGW33PEM2Q4eDjPlGi8K+QXQ+b0ucrpT9/ntMHM/wMyJggiL17wuNW4mo7dcC6FGI5wABI8GggYAmeiqFr0rHkYUcqjQJpLYaSff13fxX8o2BRfh4M86HnCqb1
D9UDu39KHlcN7i9yurunqhBRkmfHv0TBNLAVZQDhMRl1wLoUYjnAAEjwaCBgCZ6KoWvSseRhRyqNAmkthpJ9/SksgHaxWJUmGGthPi8iGxZ/WM/VJQ5ep1nWYtshQ1yI
HvDkcfoZug0a8cuoVesR6jRi6/Q7+mjbCiqWtUGmNqz+4cAuvSY/V58BDExZGMNsu27PjZTUBeQrypVjI/uWHZjz2qz8LtzUgyMcwuPyyjSaBgmuZEkASg5OzfQecgXm
kaUI6BdDB4cBakAqvDTW0nHGz7FO4O7G3479t+2InFjDThk0HSbbuy/SuJkQkbxpuNYUigRXROBTHDpltqRH4cqIJtEmvYeBjKtfeWMCbYirpY9OqzrTG3VR9UcCk3LY
nreOuqgKTuhm8gA8sOhYIVJNF6P4jjkcrSioL7yu0W60apxMwga4HaLZcUHNGSDhR2xPEdIx7xRpEQD2z8jxgeHMXvlvE9YudIhbqk5DGND/WjxPbB+zCONnzyOHdWt5
eRER9FFAT3UsTdMkQZoRTRP3f8LEUfd2o1rINGbjZ6PuMif/eUQCsS2aKhtVvj4pWKWLuou56+3z1QOZo5iLoWdyQjWL9s7MOjuGNxYddafZg8Goa19bmST21RD1oNRU
cARe1PME1f0AJ/rJQ4AKvk8VkE5SNQvAY1Mih8waGeIe8ORx+hm6DRrxy6hV6xHqNGLr9Dv6aNsKKpa1QaY2rP7hwC69Jj9XnwEMTFkYw2yjfsWuKq5lr+IihlDWJbcy
67yBrpvrBP/q4kT/GpxqJcvvygXEb8unvqp/5eSvJQqHWZVFN1C4ZdsqpdxEhvEcujfnf8LQmPdlSAnpAsgap7qo4MVa0I9vRufFLah8e6wSsevjo+Vv27W5iDVIgfdK
mgYJrmRJAEoOTs30HnIF5pGlCOgXQweHAWpAKrw01tJxxs+xTuDuxt+O/bftiJxYw04ZNB0m27sv0riZEJG8acLoA4K1iehCh5CcSvXpK43jUWd8J5mQUmZonBqVVrmE
q6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCFSTRej+I45HK0oqC+8rtFu1KeaND9mXXUdKeTmvF+ALX9Yz9UlDl6nWdZi2yFDXIge8ORx+hm6DRrxy6hV6xHq
NGLr9Dv6aNsKKpa1QaY2rP7hwC69Jj9XnwEMTFkYw2yjfsWuKq5lr+IihlDWJbcy7hn7gTaNlWV/YQOI4h3Q+sqIJtEmvYeBjKtfeWMCbYirpY9OqzrTG3VR9UcCk3LY
nreOuqgKTuhm8gA8sOhYIVJNF6P4jjkcrSioL7yu0W7WUvB2GTfY60uSRmXbl8XWqg7w03osV3q3/l2i+eboiMoo2YfC5sH4iom1/1pAsmTFxot4a4Ehzo//xgaGY7Kc
bb0ZvhE+fOZNNdn4Dk8m+97YN+iWSI0zfA+1UPUf1bJb1AyFda9cO1T5FY3kfb1ij3d9D3UXozMAstxgm1GiJ+vtgYcisHDv1lVcwx9z2M9QOrknyVnEWAL3FiNu/aIA
HCbwIb9tMK73zoatBAt0hc4zLCah9DO4zlitHEIUDba9j4b+2WyrQpbTopmuMgK6siOeRKBCBKJAzYw1Ewm/ecXGi3hrgSHOj//GBoZjspwofF+5BfqhltNQZmanSAxa
0tYsKq67owebpsuuCNaqg8oo2YfC5sH4iom1/1pAsmTFxot4a4Ehzo//xgaGY7Kc3WGp1YV48LbSwTfm6RauU0a6BDNp387rS3IzNKsmJYCTUZmc6FjBEvPzR9vujdoa
GxbfXavHOkXhfnfqHO2TKl1uKb5IoJfqM8lWLwNt4mlt2hFLlc8LQ/Ink0BJ0reaHXFUaBdcPqFXsErURCkDjOu6BmvksZPrPVnkh//9g6nwYI7d3Cz8vGNhQbTRMJPs
mgYJrmRJAEoOTs30HnIF5vrscHMSSZCejGsP4cxCmQGy4aBji6WrZpfZgoMszWEjtOjHwQlT9prK98XHltfEJuTEx8AjzXJ7P2jEV4w2xN4dcVRoF1w+oVewStREKQOM
EQNeT0ADXzgBH+YSSlEgOgq9++V7N7TaeT9yULgxf3pEx7SDuyF0S5IAc1wGiFcJTQgpui1kSkD09TMlH3otg3vZeKBTeizQs5H/wmE+OpCmhFyOO5QtzRUy/XIu75cZ
cFZfXSWvI+nGKVpcfce8gmFSpK8LoSM34kzUGWh7HETNIb0us7Sh4bhF/lTn0oGAf6MHBfOH3c4OyPtpP89+l8qIJtEmvYeBjKtfeWMCbYhNCCm6LWRKQPT1MyUfei2D
e9l4oFN6LNCzkf/CYT46kGEHVKFOdqARf8UW+wsYSNWeXNBbevXX5FoH4fMuRNQMfEEVTCEPJAt3Ywcvx85ikyeMmuho0XzM4kd2bV1UNokip4tmTuvt65r3ZpdTkk7G
wdBTD/s6LMpMggtF1i1tuLIjnkSgQgSiQM2MNRMJv3nFxot4a4Ehzo//xgaGY7KcSovp5v1Q/Ic8eGjSVSHx5A5e3wX2cTBhRDGyMBtNEsXcD8/GBBhaBgkLK12fVWpR
YVKkrwuhIzfiTNQZaHscROt1yFYHbJv4YH0chyMtePl3NhFJimsRasEAGHoikDVHyijZh8LmwfiKibX/WkCyZP7xlo3xS12ZJFxIIMx3LG1UuZ/4YywHdYLj1Mr7wE2B
FPKEArEApczWfGkIJVSlKVvUDIV1r1w7VPkVjeR9vWKzdLcjZ73/w5PJl7jvXccDcWEpqyjo1PwmJLaNLN6gLrscyheMGBf297+1s5w5SCNb1AyFda9cO1T5FY3kfb1i
s3S3I2e9/8OTyZe4713HA8hCHPCheslXMUMukcrCvmdwVl9dJa8j6cYpWlx9x7yCYVKkrwuhIzfiTNQZaHscROMAzSNJL8aIj+Eq9fbvyKhFYDecDkBvgZn+lEGu6OLC
3A/PxgQYWgYJCytdn1VqUWFSpK8LoSM34kzUGWh7HETjAM0jSS/GiI/hKvX278ioIzFiyh2ud9mJ6B0USgXROdwPz8YEGFoGCQsrXZ9ValFhUqSvC6EjN+JM1BloexxE
bNjANMVb7cV9YcDBKDW+lbpGPjWm9Td21xrd4STsflq2glUm3FiRKNbzicOYw7arJSOqmHfq4/01r8uJCDDAR4Z3I1Hd4lx0DqHs9MdjJLcgGdqO+/GFWgXX9XRPVwAt
LdkpiGwU3wtS3/dM1DZIa67sFiZbfPhgZz4WiRR+3rufH7NZdl667JFqk7Zr0zkHnlzQW3r11+RaB+HzLkTUDHxBFUwhDyQLd2MHL8fOYpMZsQoB0W27O2vZiV/nWMrN
LpGT4S2HJ3+2SMQPpJKnlsqIJtEmvYeBjKtfeWMCbYhb1AyFda9cO1T5FY3kfb1ilgMndTOBrI/iKs+CeopHirNP2G0yANdsWVaDp2Z2R7PcD8/GBBhaBgkLK12fVWpR
YVKkrwuhIzfiTNQZaHscRBGFAWydaXmDzELTQaM8R4dtvRm+ET585k012fgOTyb73tg36JZIjTN8D7VQ9R/VslvUDIV1r1w7VPkVjeR9vWJapcrzqqNjrSgCYjRfFbYL
RjFOkyrR6l2IrnxQdobYvN8ctBV9iAOJmsnxuiIIJOaJADAh8iZTFIsekhFmhwlEGbEKAdFtuztr2Ylf51jKzajDi9b69o0VLqf/U39KFcIg4bhbVoVNR8l5+tmh9qcW
czOnC534/bgvwa0RypMZvfOIswZFqGrG+LaLw/voDkmo6zXr246msXmwuQz2kM5/KFRyCjG0vmqbFWeswnv7pnxBFUwhDyQLd2MHL8fOYpMZsQoB0W27O2vZiV/nWMrN
Nvyh1cyC5iBA3hP16lmmOq2WPl3UpB+JWOqJkkljU1dzM6cLnfj9uC/BrRHKkxm984izBkWoasb4tovD++gOSVToyBCmnPW8//wUJUFQ8YM21edd5XN/3hBGKeSz/jQR
azL/a65HSi89prYJSVrX1EHdgbK+zP160x6kSbSiy3U3ffspGPN7YRugkwnIGKOfwdBTD/s6LMpMggtF1i1tuDR/oh53SoJMAsUaIXmxsb/+8ZaN8UtdmSRcSCDMdyxt
Sovp5v1Q/Ic8eGjSVSHx5BWdne0500DZrSfKeQkY3ohwVl9dJa8j6cYpWlx9x7yCYVKkrwuhIzfiTNQZaHscRBGFAWydaXmDzELTQaM8R4dtMMuN226dJ/btcAQiufha
71BFeVsA7K2EsdtazfFyjXMzpwud+P24L8GtEcqTGb3ziLMGRahqxvi2i8P76A5JCk1+Y6Vxga5grwEePdkXD+I4tWUfFltSHSTAAl2qG+DR5ShRIl94UvBsC1M5FJnJ
Ii5k0S84V6ZS8qOAXMN5VTqYcAEy7WgOQtBKCKCtVfTFiupUpkrgBtPqTrrf311BwnhpVTvwwoJr/ftGExDiEyo0kjYRofXmlqdnWqJ/5wnATnCkUjaz3KNWBeacD8Ff
LiBtMH5vpNjtuqg0H7krGcqIJtEmvYeBjKtfeWMCbYhTpuA7aHOlUzvSIMDFGxtbwMjiTqX8rGSnOBxzD3sQf+VhExDcSrj8oi54pE37vXvsVU3OE2J7ycTS0x0spYZs
5yIM9OdllrMKvacu7WJvC+FzcmBY5eLreHNcckBJcsB9HADgIijAhu8JM+btDKhY7DFhx+bklAnVUt7ltfN6fcAKXX63Ck7+j7kx6Xx7Kx3v2ucU1EoJHGNjR/0HF0Pl
tKLjYKJs4z7+MQ8Y2jdbI7CQSjbG/kVqerVxs63q3zltHSTLpes4HhzMSie4S5GK0LbikoFrpXimYp3cTP3RoEq2qUlKZVFpnMWiTRCiuFsq/NG/OQFjdXnCdVe4ITZs
3SqR9IuGx/LgCWP6V834yS3tyb8ZAl+jJmZKxy7RPuaWR+JWi6+ySV+A7JH99vIeVSHn0RFLrXTPvg8oVw9CKh86rjKkb8nghKApTXhTeQw1rA1AuL2OCkuBxawLwaB2
bdoRS5XPC0PyJ5NASdK3muciDPTnZZazCr2nLu1ibwvhc3JgWOXi63hzXHJASXLAcDvwSK1J0kCMnNPZN5GdNxk2YQ3HQLPxuqXw8Ts+lmEEz7OH7NQB8S0bGD5jOdV7
Q/wlCVvlysRgS2xZTi6sZKkEofYL2Vt8CT+Zq2w7U0Qo3uTf/NrlvMExTlVbTVNWhtI/Vu8MJaYwqhb4WZAsFDzf7f/Omwvyit2r6CcF7b9Mk7aOs58AkAS7w4D7A0lz
XZkceqaa2kAP91EEvYntBo4R8zJhe3kc+ZAXe6nIBLaPAr/vhV7nA9dhRR9fGysNgSEUBihJp7fQjaAWxz1C8ks1iy6vPBLkgjJzW5M4znG/lQs6W3xAGhV+3WI/bZhm
lyTeHUSjIS6t5D6V5b5NA8qIJtEmvYeBjKtfeWMCbYhTpuA7aHOlUzvSIMDFGxtbwMjiTqX8rGSnOBxzD3sQf+FB8sW+I8iitd1pElnWIAXkxMfAI81yez9oxFeMNsTe
5yIM9OdllrMKvacu7WJvCzgDP5Y9snkQBlO1dgjIvCbtyUsOJD3CS85a7SzIsCE7y+/KBcRvy6e+qn/l5K8lCkMN4PSPcUN5UaU3Wq2lq1o69dBpGbv2JcIFeS3Vw+wm
7jIn/3lEArEtmiobVb4+KYqsZh7Kpflbox+GsqFkva9tHSTLpes4HhzMSie4S5GK+ylDZ1EWKgRAYoWvuybFc49msKNMg75D69bo/5X2YmpVIefREUutdM++DyhXD0Iq
HzquMqRvyeCEoClNeFN5DB+fhGev3eQ0ZF6HTotF90SaBgmuZEkASg5OzfQecgXmBM+zh+zUAfEtGxg+YznVe5OfNef3l5VwJTsTaOXPGaRh4YAPvw4jNAzwO9MVn5FF
yP5Pk/x2LpeJ54DVgmXd+o4R8zJhe3kc+ZAXe6nIBLZ9/xdmvPug1WVPG0IOD2Y9R2xPEdIx7xRpEQD2z8jxgUs1iy6vPBLkgjJzW5M4znG/lQs6W3xAGhV+3WI/bZhm
ab/PxyVuVEKcIsDBWZ/+Ebr/d6zTt+cL7zyOVXqI7NBErqrRWguLLMviEzmaZhjHcZWy5lc6uib61r2GeIexqwWmsXj2ah0jEAWK/qPR0lVEx7SDuyF0S5IAc1wGiFcJ
U6bgO2hzpVM70iDAxRsbW7dh9n5X4tHBSzXSq5xqBmgepRzzNXw7fnFtOimhdQxAR2xPEdIx7xRpEQD2z8jxgUs1iy6vPBLkgjJzW5M4znG/lQs6W3xAGhV+3WI/bZhm
w3/rZKv9d+OuO3B8J1riRdwPz8YEGFoGCQsrXZ9ValFErqrRWguLLMviEzmaZhjHytXRGI4e4cssMYMDqVjjo721jSWOnkx+HKg0SkmdrkBVTFcJNWYysVpHtG7kevqG
wApdfrcKTv6PuTHpfHsrHf6yINodZ9ljy98l1wVzcke0ouNgomzjPv4xDxjaN1sjsJBKNsb+RWp6tXGzrerfOW0dJMul6zgeHMxKJ7hLkYrO3JFtVLGaChp2LkqCyXXd
cFZfXSWvI+nGKVpcfce8gkSuqtFaC4ssy+ITOZpmGMfK1dEYjh7hyywxgwOpWOOjko6r2p24EFGxD7vAKUjai8vvygXEb8unvqp/5eSvJQpDDeD0j3FDeVGlN1qtpata
D8eYg45tRjpskhNpianu2ZDdT2rcUC5+gEQ/BhhH+/XmYZrzgb/FN7VovGbra5Y8dwqEgAVC1UcVDpdJHnW+s3c2EUmKaxFqwQAYeiKQNUe2t9evRLSI+bp2ZNET2bku
v+TnZzKxiZGKq6R0TUkR/721jSWOnkx+HKg0SkmdrkCWzti7uOPipdwPmbYudIKX7Y9sIRX18HkUh64DK0pygcBpNhSiZKTA4NBZrqrG3qe6+9x0TU1U+1qDZgR5SMhe
0SauVx/M+eatLe4uvcRhH/3KXbzzWgjRzrCGczMJsyC6+9x0TU1U+1qDZgR5SMhe0SauVx/M+eatLe4uvcRhH7Xs2f2p3xb4RL5ROxZZrvyLBQsXlg7+6jxSUEou9ylZ
MXt8O19o3CUowtMPmKGJwry/m84Va5pyOrCI/wUoGcQdDnDV4VvQlhOsqttR41jmMZ+AW6CuIynWQ9SXnhj7FdWuxkcD/ZAbnV2Rgyhkxkog4bhbVoVNR8l5+tmh9qcW
I7uonJSw1YQ9XLGHuIjY/Lfp4yM5X+VTS7AahqhbMVcLoDmqlfjNoP1jM/eiYw7SuqNtEGSQNT+HsQnmdwxXo4eoEwwnGntXI518AVMjLUGpBKH2C9lbfAk/matsO1NE
inwS07r9Hh4LSMCzBBGrhFxSXg0jjJFHnwAHXIi05UmrRU10XbAqFT2AH2j1tdBx/ozHgkCqtaWGn4lSW4utgFf9ivgvLvDD4xtWEufw+3meR1xl3agwcJpXSmQCFK2o
ugpN6ETPpj4hVLqyDp2LJdEmrlcfzPnmrS3uLr3EYR/kro7wCXolmzMdWSYg110A3A/PxgQYWgYJCytdn1VqUX9ngNZkSSSWWO+ecUbmphEl6GO9M5RqtUbeIXUQHfzg
Vwx+DswoS4b26pi174TNQ22ggoMsjkBwPrhRP9KkgGeDMJXs+7m8IRpdzfVUHKFdSL/qdzYJN6rMuUFYw6VK043r3bzM7n2Lz04uEcMWtTJ/Z4DWZEkklljvnnFG5qYR
qqIunUMe9ROKyqM2j9gmVw9599uYJgDHN/4piCTz92pWRzWnO/TKWSQyMcBOkpeKeeaofWixv60vDrnh9shfQ4gjr6lkYvuplshLA+RkwZ0jIIQGdUUiQMU1qqA+UPWj
7Y9sIRX18HkUh64DK0pygSZYkpcs9Wu3TUJa4u/Fwqnh1ykjBMmUP982+jC0BNalI7uonJSw1YQ9XLGHuIjY/Cg+vrW9xFhmrvHetGFVZI5iAgN0CP6xujLlgB0AqzAf
vNDlLdqzDjTe04NbDuj/jAwccNaCslQ5EBZwjXODP+VSy+xuhbRr6RJiUfsLMbawcOp3fPg4o+gTUr50Ls0akTF7fDtfaNwlKMLTD5ihicJ/99r9aZ1jirkQAtLk4G0P
L7gortYATjPI6kElQO4NgMFM0vXM/N3TdgS3RJDSZVdcUl4NI4yRR58AB1yItOVJTROqekArkTbYUess7SWJF+aNhkZM+nHl8eQMfXZp5MYFTNf+juK880vz8jdPp0Nw
duSPecRWy0uUaTsnHPOmI6I7OeKYxx/mcdSlwpZxrN9HEQilmuoWTZ/gFaV/8dnmv+TnZzKxiZGKq6R0TUkR/w/JnRMsH3L9hN1hQhzbvCedrcYb6SYtCMfymE/qt9vg
jbbJiPB6yi6fj23v71W2d5BkHTTjrmlHEbBFt1B8sk+Q3U9q3FAufoBEPwYYR/v15mGa84G/xTe1aLxm62uWPKj7lx6rGZXI0sYP7il6kxR3NhFJimsRasEAGHoikDVH
trfXr0S0iPm6dmTRE9m5LqudKnSHFFnogOY+sKZafFq9tY0ljp5MfhyoNEpJna5Als7Yu7jj4qXcD5m2LnSCl09YKziAbWW1a7gmqZ9YK9fAaTYUomSkwODQWa6qxt6n
uvvcdE1NVPtag2YEeUjIXk/qWBDUi0LpH7WXTM9ERAD9yl2881oI0c6whnMzCbMguvvcdE1NVPtag2YEeUjIXk/qWBDUi0LpH7WXTM9ERAC17Nn9qd8W+ES+UTsWWa78
iwULF5YO/uo8UlBKLvcpWc9QSEevqjIAxGIz+nluXuS8v5vOFWuacjqwiP8FKBnEHQ5w1eFb0JYTrKrbUeNY5tR0HBnMiDPcNOq8a/ppOf7VrsZHA/2QG51dkYMoZMZK
IOG4W1aFTUfJefrZofanFiO7qJyUsNWEPVyxh7iI2PyUjHqki5pNChElyswYRDBRC6A5qpX4zaD9YzP3omMO0rqjbRBkkDU/h7EJ5ncMV6PHbRXHf5Zf9hu5ampD0G3K
qQSh9gvZW3wJP5mrbDtTRIp8EtO6/R4eC0jAswQRq4QtAs4dxocDQJETu1P6IB4Qq0VNdF2wKhU9gB9o9bXQcf6Mx4JAqrWlhp+JUluLrYD2QhwfgwS8bgrmqC8l4rjz
nkdcZd2oMHCaV0pkAhStqLoKTehEz6Y+IVS6sg6diyVP6lgQ1ItC6R+1l0zPREQA5K6O8Al6JZszHVkmINddANwPz8YEGFoGCQsrXZ9ValEwx/VUQ50AFR1219X1QbGW
JehjvTOUarVG3iF1EB384FcMfg7MKEuG9uqYte+EzUNtoIKDLI5AcD64UT/SpIBnltH1GOWSY8vyZ2v6qDEC6ki/6nc2CTeqzLlBWMOlStON6928zO59i89OLhHDFrUy
MMf1VEOdABUddtfV9UGxlqqiLp1DHvUTisqjNo/YJlcPeffbmCYAxzf+KYgk8/dqVkc1pzv0ylkkMjHATpKXiuQN8SM7sNvT7AIVDrzE/OWII6+pZGL7qZbISwPkZMGd
IyCEBnVFIkDFNaqgPlD1o09YKziAbWW1a7gmqZ9YK9cmWJKXLPVrt01CWuLvxcKp4dcpIwTJlD/fNvowtATWpSO7qJyUsNWEPVyxh7iI2Pw5fxZkIrbDoJAnTMlKAokj
YgIDdAj+sboy5YAdAKswH7zQ5S3asw403tODWw7o/4w2UOtyVY2zRYHSzPRD/6pNUsvsboW0a+kSYlH7CzG2sHDqd3z4OKPoE1K+dC7NGpHPUEhHr6oyAMRiM/p5bl7k
f/fa/WmdY4q5EALS5OBtDy+4KK7WAE4zyOpBJUDuDYDBTNL1zPzd03YEt0SQ0mVXLQLOHcaHA0CRE7tT+iAeEE0TqnpAK5E22FHrLO0liRfmjYZGTPpx5fHkDH12aeTG
mjLgQBgRAdsXjhpzErIo83bkj3nEVstLlGk7JxzzpiOiOznimMcf5nHUpcKWcazfRxEIpZrqFk2f4BWlf/HZ5qudKnSHFFnogOY+sKZafFoPyZ0TLB9y/YTdYUIc27wn
na3GG+kmLQjH8phP6rfb4Fhn7rca2mmehrW9BM2crGyQZB00465pRxGwRbdQfLJPkN1PatxQLn6ARD8GGEf79eZhmvOBv8U3tWi8ZutrljyDXevbED+b9FmV7bUbifGo
KkHTYLZ3eFVgR6Fcq8b8rPGLxF3AJyF4IFHPHXeCOOzJHfFUxnZqhf8lD2tmOBPQykpcuO+kuOTpVU/Mw09qmlzXcQDkLRVCJX4hpHNAmE/Z7Po0klzcD/dAYZKPLkIE
ju9N5hABfYn5G1t2EH3j8br/d6zTt+cL7zyOVXqI7NAOQSonnyZJLWKpUupgzNe6lXpWb0YR1W5aCpYrA5R2NzPEOW9l12ScTCtyYVqrwQptoIKDLI5AcD64UT/SpIBn
2ez6NJJc3A/3QGGSjy5CBCMxYsodrnfZiegdFEoF0TncD8/GBBhaBgkLK12fVWpRDkEqJ58mSS1iqVLqYMzXuknp0plYD8pJgdzr0HbVhiL5ddCSBTIo08r9EQ6D3+L/
ATS3T+Cof5iHKzJ3RnS+xIZ3I1Hd4lx0DqHs9MdjJLc1iIeteFOShEHQjXD4OIR8uqNtEGSQNT+HsQnmdwxXo1xpJLwul+Db3Lz80RyBWe+NosrGEQJ5Cb48Pf08Kq+D
gBUXChQW4jk9V/40iULYjeFLm5ztLvzL/b99qlUz+rsJzr8LICsgEXo7XZ6gx7H4R2xPEdIx7xRpEQD2z8jxgRpDvz1GnL3RsFSurpv0r0c6mHABMu1oDkLQSgigrVX0
sgU2Ffh8TSIauBvH6H0iJYAVFwoUFuI5PVf+NIlC2I3hS5uc7S78y/2/fapVM/q7JvFoETu3I22n+nfHj9Pi6cpKXLjvpLjk6VVPzMNPappc13EA5C0VQiV+IaRzQJhP
yFXqq2r2vPWuUQD83fekn2OXB3SHHmvfVd4INin5Uz/mjYZGTPpx5fHkDH12aeTGuzC29FwvVlIqyy+etodH/GKxR0NPLVsXgBJz1rGYsIcjuAZHMUApoIovmVYcI3M2
EcfsZ5yjd7gxtzIsHi9eQfrHJfoXZW8Wmu3XKOSA+fNED14nSJj8XohTrlHzGLyXt4tonZ/uPsgF1gg/bcH8qzReh7fs+XhBiyhXHAVUDudAt9w3BZXKqVM8UkrHqlw5
eeZQv7xEuJVV4PgeIXMOFuCsCD3UlWynLeS4fDBjEsbhS5uc7S78y/2/fapVM/q7u27PjZTUBeQrypVjI/uWHfbisAgDD+i6KGoKIEb6/jr+jMeCQKq1pYafiVJbi62A
gB2OQzVk0Mc5OLbZA75WeApNfmOlcYGuYK8BHj3ZFw/ozUUIz49GVJ0hNgja8njoRm8zRLvUyoKOl2L0/9WwCpxxg0mo9YQFRpeuQs9iANQip4tmTuvt65r3ZpdTkk7G
kOoC/wtscouWuE1hL3U6XcvvygXEb8unvqp/5eSvJQpkXDcEO7m+RbsSCxdjNRjKPj2LnFcqkwkTtXk+hSznClIFH3NJUTH+Y4Nca0Q1uaTKiCbRJr2HgYyrX3ljAm2I
U6bgO2hzpVM70iDAxRsbWz2UHhRP5OuAUuUz9JhC5sA6CQRBYHFStD0jXNXIUPR5hN4LSGBgzYA3AaqvHjYDIxUbvSNA0StMlLdEhfuPecBkQqy2K9YjZeCH1DEP2Kr+
7lBM0H+FFO4L4RIVIyvinVGfKvss99kkAFlBAcwKnwbsMWHH5uSUCdVS3uW183p9CJwL3yI2oXIWE/vNov5Btzc/GciEbh6eNcCkL+wsnNs9tmpE+FKXC/CzIhQGpn/s
bdoRS5XPC0PyJ5NASdK3muciDPTnZZazCr2nLu1ibwvPp7rkEuLbH99Gdc/bGq8WuNWuAFPd6zcTryUW1QWgkkdsTxHSMe8UaREA9s/I8YFLNYsurzwS5IIyc1uTOM5x
f+FNuaQkD4OekxUsPIitdExiw3h+FQrhLsbYoA7dwOJoT4BhFhMTECGmG8MrJQmiyijZh8LmwfiKibX/WkCyZOAIDQ7985dEFe+Zy9ggHRGvZIKsej/gpWjbtnYAnMeu
LW53280uqMkncBzWtNEdFI3r3bzM7n2Lz04uEcMWtTJErqrRWguLLMviEzmaZhjHknchx1kkk/tqGcwEsZtJGSKni2ZO6+3rmvdml1OSTsbjgUjTDbKrphgFbjkbbrv5
3Y+e4YTMDjyZicr+JJtWH2RcNwQ7ub5FuxILF2M1GMo+PYucVyqTCRO1eT6FLOcKnx+zWXZeuuyRapO2a9M5B55c0Ft69dfkWgfh8y5E1AxLNYsurzwS5IIyc1uTOM5x
f+FNuaQkD4OekxUsPIitdJWnE5sPFEBDdKjcB2LOiu4GXuPEAQQoaIXDIIizxe1N5MTHwCPNcns/aMRXjDbE3uciDPTnZZazCr2nLu1ibwvPp7rkEuLbH99Gdc/bGq8W
j+g69/0HrnvS5drhxr3rKtt4mowQsID/3OY/vgLUyGvrsK1wupmEpoCynz/bdPSgVnVeAHPGGg55wUkV9hUNHhmy34mLa2bbiuoyyUvtdUEpSJDo17mStAxRbrOW9kGT
3A/PxgQYWgYJCytdn1VqUUSuqtFaC4ssy+ITOZpmGMcJ8imp3qNzXT8cupIVdfwPYsNPoYNN2ME5ZQLfmFU1kbDPrCzgt8ho6MTxoAaPvYkq/NG/OQFjdXnCdVe4ITZs
KUQ4MOY8TOL4inlOOB2rQ/SSgYmgSh+5ss2Q5xP4yzEFprF49modIxAFiv6j0dJVRMe0g7shdEuSAHNcBohXCVOm4Dtoc6VTO9IgwMUbG1s9lB4UT+TrgFLlM/SYQubA
qlfy4aAp+MS9Ffap7uT2D3lzX4nnp7uQuAbOfn4FdY+AFRcKFBbiOT1X/jSJQtiNSW9NF6CKBuHLdrfZ8dEq9qQgLfaVW9wip5l5kSqsCglm5V0F528oOueXKR/h0AsO
IUj20Fdxg5KMSTkjetcNp2Lw8EONRTiCKVwTP1lZJpWuLO+vk5M9FpJrEpM5cq/x8a0W7Lf5Brxz9yEwEbS+Xc3USAdZPZAbq6W3+7igQEcxLFNhjd3n4e2W74alQGlS
SW9NF6CKBuHLdrfZ8dEq9qQgLfaVW9wip5l5kSqsCgkt3JXg+oQT4WfTOhh+TUFE82H2XK6oLfhprqp8qkgIXsoo2YfC5sH4iom1/1pAsmTgCA0O/fOXRBXvmcvYIB0R
6kwi3E9EpahpqXhQR7C9pgxcteSq/534zfTmJqwjBJJp9x/TVikdNR+F1KSEHESYyP5Pk/x2LpeJ54DVgmXd+taPD5cDIrRUHT9uMwCaPT8MBF4R0XjuPq/WQPKOD54G
7PqI7CXnHqIxvghz97+oyrSi42CibOM+/jEPGNo3WyOwkEo2xv5Fanq1cbOt6t85ZEKstivWI2Xgh9QxD9iq/hgYoVQenuAY6boPS3QxABRSd65LUpRkl0bUQsIEVZ15
K3jLMlHAzBu0+n689gXkESo0kjYRofXmlqdnWqJ/5wmiSJm8zvSwzWRrL/xDAPy7TjvgjRuEuQ746kLwRD9W7n+jBwXzh93ODsj7aT/PfpfKiCbRJr2HgYyrX3ljAm2I
U6bgO2hzpVM70iDAxRsbWz2UHhRP5OuAUuUz9JhC5sA2YCEAUJAJ4riSwfLUO7S5QyP2gpZ0DxQjDsF3O2Dj+eaNhkZM+nHl8eQMfXZp5MZTpuA7aHOlUzvSIMDFGxtb
PZQeFE/k64BS5TP0mELmwDZgIQBQkAniuJLB8tQ7tLlUiPd5uLma4kbEkN8Fk9hfRroEM2nfzutLcjM0qyYlgCo0kjYRofXmlqdnWqJ/5wmiSJm8zvSwzWRrL/xDAPy7
TjvgjRuEuQ746kLwRD9W7iOP8EqFNrjvBiFSQu3pux0qQdNgtnd4VWBHoVyrxvysDlnCS4SR+JHwqj0zdMRHHY64hFGigmzSxv33v/XbSZVPHnev8P3bhs2CTtb5zHxu
3tg36JZIjTN8D7VQ9R/VslUh59ERS610z74PKFcPQioAWLNDlpkRPs5NxIYIWFq5tueDTG02eV391IQuObuPqeCjrbOm6qMfi3YL8s7iuMysOBxp7Ockz5a1S2udZx3c
c/Rfo55o5WKosjshnvyoGrSi42CibOM+/jEPGNo3WyOwkEo2xv5Fanq1cbOt6t85jriEUaKCbNLG/fe/9dtJlTGj7+XAnMwn4wabkWHmJR9sQlaQqXt+jNMreIPOEvi0
5yIM9OdllrMKvacu7WJvC6V/H4LC56YqZpLvuF/eEFcA9yhQhu59m1d87351rsN2QbV5de0XGq0UmAe1pUQao4v+z/HuxEsny8q6WG6duGJ0ZGpvDrNuIbRodkQ0fY3T
gSEUBihJp7fQjaAWxz1C8ks1iy6vPBLkgjJzW5M4znGfHXC/bRo475erqvIc+MXIsncU+aExtBTLyp5QO8IFRDEsU2GN3efh7ZbvhqVAaVJJb00XoIoG4ct2t9nx0Sr2
8LPtX/h5vx0qDARnQ5y4YH6rYwpGcr4E2Uxdh0mXvMZo2MBLOkM3JW1YJuk/IZ/C1I7avMtgryDQY3vGHp32rCJPeXyL0y74S5IIGKY40dsKDLQ0qQCNovUuexI/JyB5
KjSSNhGh9eaWp2daon/nCQJYhHTDzXpYCQgrDr5yyn/nfDefwRynsaDsu10PNKpBuvvcdE1NVPtag2YEeUjIXklvTRegigbhy3a32fHRKvZstsODlAN4xuWudS/1fj8c
fxcLnQylypxZnRLmA93hsLCQSjbG/kVqerVxs63q3zmOuIRRooJs0sb997/120mVI1lRNBBQBj8jmFRYHkqm5MqIJtEmvYeBjKtfeWMCbYhTpuA7aHOlUzvSIMDFGxtb
NUDItG+ZqffIknp9m51ls+1YFhsNROIEaScFJi78lNjR5ShRIl94UvBsC1M5FJnJ/pSHMoFnljdB86Srl3rzZcrgGNxqvvFtJ052TO4R6CGtlj5d1KQfiVjqiZJJY1NX
YvDwQ41FOIIpXBM/WVkmlWx74GoJyO9XEjmz77yLuOHqV1iAeuzw8YITAXTA3PtBse4GYyN9ckYCqCE6sYDPY0lvTRegigbhy3a32fHRKvYeZW4kweDHZcUMhK5Syr35
rjxSPg1ZlLi9t52JVLAtPzoDFfsfu+puZMausS9a02dTBmoWuZy0yJa+iGXEQZ9F78Auu1DaQMN9BsKFcqx02YAVFwoUFuI5PVf+NIlC2I1Jb00XoIoG4ct2t9nx0Sr2
2b+x9aEsLyVZxoyEHaHOI5DdT2rcUC5+gEQ/BhhH+/UEAryO2LIZOMoPRLzF2cA7UwZqFrmctMiWvohlxEGfRT8WQtx6+vv4QHa64Rc6fdrkxMfAI81yez9oxFeMNsTe
5yIM9OdllrMKvacu7WJvC0uTW9iaNmMmQsByC9X0cbjKSly476S45OlVT8zDT2qaXZkceqaa2kAP91EEvYntBvD1Ga78B8bdjzVYgNp1r9oQ6r73QFA9lP6LzuyQbeaM
3rdgMwHcs5xHKxXHDvdw0Cr80b85AWN1ecJ1V7ghNmxTBmoWuZy0yJa+iGXEQZ9FHLeDk6/GCYhZxJmOCcmt7JDdT2rcUC5+gEQ/BhhH+/UEAryO2LIZOMoPRLzF2cA7
UwZqFrmctMiWvohlxEGfRYNu8YFh4wXpK2aWoQdRgobkxMfAI81yez9oxFeMNsTe5yIM9OdllrMKvacu7WJvC7bo/wrSjyWOhttmIyJkJfkqH3dTFVR6f6LDt5uHh4fR
nOQLCZocypSRUWGe4rodS/D1Ga78B8bdjzVYgNp1r9rvwkTn/akm2KdlO0MM8ZUZuv93rNO35wvvPI5Veojs0ESuqtFaC4ssy+ITOZpmGMf/MSXUl6t7oHPv5/ugHoQJ
3rdgMwHcs5xHKxXHDvdw0Cr80b85AWN1ecJ1V7ghNmxTBmoWuZy0yJa+iGXEQZ9FDZu+0Znje7HHnXs/92gC84AVFwoUFuI5PVf+NIlC2I1Jb00XoIoG4ct2t9nx0Sr2
TMoD8iMvzYnGwNLO0hZoy5DdT2rcUC5+gEQ/BhhH+/UEAryO2LIZOMoPRLzF2cA73SqR9IuGx/LgCWP6V834yRet+511oPw4YwHi7U6syAGyBTYV+HxNIhq4G8fofSIl
gBUXChQW4jk9V/40iULYjUlvTRegigbhy3a32fHRKva8l1x2c7AW+LhyzgcZORhlniiOPBly3YabwwUaQBlMF4vKvqUAxMn1Yx/4GLU9PJU6AxX7H7vqbmTGrrEvWtNn
3SqR9IuGx/LgCWP6V834yRet+511oPw4YwHi7U6syAEuY9X2H99YZ4xCbIWifn0P/ozHgkCqtaWGn4lSW4utgATPs4fs1AHxLRsYPmM51XtHtWffV/a/nQDDLRn5KJOU
026xh42rjzDD76d9+qdlGCc9TI8VVfxwqk77JJv5rchVIefREUutdM++DyhXD0IqHzquMqRvyeCEoClNeFN5DKu3dUBInu0gQUvkuP2C6FEA9yhQhu59m1d87351rsN2
QbV5de0XGq0UmAe1pUQao0MN4PSPcUN5UaU3Wq2lq1ryJGO+rSjRl3AeuzqsNGyFPllFepfXs/8ZMpjlGlmZOZB/keYmgETpbFXygYEtO2pTpuA7aHOlUzvSIMDFGxtb
wMjiTqX8rGSnOBxzD3sQfzCejnA56ghRjRV/nsnFm0xHNO0nIC9h9Zu+2bLSDeYEXZkceqaa2kAP91EEvYntBo4R8zJhe3kc+ZAXe6nIBLbWRIdbCnvBu7/omxlfEapv
n/OJhfwq3pKHya662RAmnc0sErjYpIovT97sYzYP+aVErqrRWguLLMviEzmaZhjHmYtJ4KB8mZWY+vKHNLPrqzPmDsnDXYytbRo+9Wg9X/C0ouNgomzjPv4xDxjaN1sj
sJBKNsb+RWp6tXGzrerfOW0dJMul6zgeHMxKJ7hLkYrHUFPVUrZY2j800MxyjiV0RH0LDhg9AvVFt2FBdOgOwmxCVpCpe36M0yt4g84S+LTnIgz052WWswq9py7tYm8L
4XNyYFjl4ut4c1xyQElywNFSwc827bzg4ogEJAZ5bVdJYySJWlq+qXWZJR8Pwqb0YvDwQ41FOIIpXBM/WVkmlcWLmIJFAjV9f1zyAzuGJEaRhYrmuGDgXzhGnrKLCFZb
3bElob40YEeoOIrZkJJTRNHlKFEiX3hS8GwLUzkUmcnACl1+twpO/o+5Mel8eysdeIRzXRNIEzQvj18azTN0Un5x5Hju45+Y8YhrltviaMriHj0rTxoZ6bRub8ATr+vm
SzWLLq88EuSCMnNbkzjOcb+VCzpbfEAaFX7dYj9tmGY6TnrhdQHpMIOPU/Sy6mE71C51JjoKkyc5KzmyN6YS6MqIJtEmvYeBjKtfeWMCbYhTpuA7aHOlUzvSIMDFGxtb
wMjiTqX8rGSnOBxzD3sQf5JMpxiOh+8fKvqp/YZ20Se1yLJ7skafgoY9fv5GjxIp4KwIPdSVbKct5Lh8MGMSxklvTRegigbhy3a32fHRKva8l1x2c7AW+LhyzgcZORhl
KJO4qf0qxCuCo61ne2pkuYzFRbWe9VSPlSxPCCUjDSIo3uTf/NrlvMExTlVbTVNWhtI/Vu8MJaYwqhb4WZAsFNJuCqPrUf8pcF7jSNahz7E4UaIEWNCj7S+p193vLyVc
Ihj/LGxdJ45k+/9siPK5Kks1iy6vPBLkgjJzW5M4znG/lQs6W3xAGhV+3WI/bZhmOk564XUB6TCDj1P0suphO46/mEQVYVRs+0G13CRGeBdYMn5zIFKlu8KVM7ogQh3l
VSHn0RFLrXTPvg8oVw9CKh86rjKkb8nghKApTXhTeQyrt3VASJ7tIEFL5Lj9guhRRIZBDtKsYloU8YESeY/0u+bbKrA+OU0N2fHXzFVl55YEz7OH7NQB8S0bGD5jOdV7
R7Vn31f2v50Awy0Z+SiTlH9G/Db16Tv/FloNN6p52mltEJmpG8XpOInf8N0bFMDisiOeRKBCBKJAzYw1Ewm/eX/hpoqEoKzZUrmj3ABtLTAAbbJrcyIIh/rwFzpZ6ELA
12k8ILn/c/0ftwlMXujDAADdEWXiSennOooQrnArRC0q/NG/OQFjdXnCdVe4ITZs3SqR9IuGx/LgCWP6V834yRet+511oPw4YwHi7U6syAF6DY9JhgxNjgdM3yLHhtA/
OUMAvypklNcCZAuAP+GyhlUh59ERS610z74PKFcPQiofOq4ypG/J4ISgKU14U3kMq7d1QEie7SBBS+S4/YLoUcg4MDBdKg70Fkbl9DYW5PxsQlaQqXt+jNMreIPOEvi0
5yIM9OdllrMKvacu7WJvC+FzcmBY5eLreHNcckBJcsDXIXTh1P36fmasYOeA+PEE2ymCIj50nV+KKXGQqYHwMLMisVzkHDO/pw0MifpxxA2G0j9W7wwlpjCqFvhZkCwU
0m4Ko+tR/ylwXuNI1qHPsZBkHTTjrmlHEbBFt1B8sk821edd5XN/3hBGKeSz/jQRBAK8jtiyGTjKD0S8xdnAO90qkfSLhsfy4Alj+lfN+MkXrfuddaD8OGMB4u1OrMgB
jUqnkDiHTdpFYQ+nxDE8OcJ4aVU78MKCa/37RhMQ4hMqNJI2EaH15panZ1qif+cJwE5wpFI2s9yjVgXmnA/BX0qxoqsLOMoQSNvg8VtjYmVp9x/TVikdNR+F1KSEHESY
yP5Pk/x2LpeJ54DVgmXd+o4R8zJhe3kc+ZAXe6nIBLYaOIIwbET4mFvje7qXrLb1tueDTG02eV391IQuObuPqVxqZMTn2+1VyHC6Vqpkh8EEz7OH7NQB8S0bGD5jOdV7
4qJHZaPNRMG+vI8+0H8+Uj3xWYL512o77bpwS0FDi51PFZBOUjULwGNTIofMGhniHvDkcfoZug0a8cuoVesR6n/hpoqEoKzZUrmj3ABtLTDkqVWqT2053kVGjS/SxRXs
bgc+MsBpLtQlVaqRiWoceq2WPl3UpB+JWOqJkkljU1di8PBDjUU4gilcEz9ZWSaVxYuYgkUCNX1/XPIDO4YkRhbeHKmKCqZxK1THO//bT+0zVcqab8gi51poCtNsbmMS
yogm0Sa9h4GMq195YwJtiFOm4Dtoc6VTO9IgwMUbG1vFKVePxJDExXR4y3mbCRQIZfNlJfMc1ur/IAYmW6OqNwYizLDg+LMiXH0jd3Idj2KKrGYeyqX5W6MfhrKhZL2v
bR0ky6XrOB4czEonuEuRivsN01MGi4gPJ37SHmkgq8oHnV1nitbzy7fmSHZPA4NGIH5X9dK/iTcqUl+BnsmuNVOm4Dtoc6VTO9IgwMUbG1vFKVePxJDExXR4y3mbCRQI
6m3l9gWBcaEL+P3e4J8wcex6uK8CWlKgT7Q8yInfRnjL78oFxG/Lp76qf+XkryUKQw3g9I9xQ3lRpTdaraWrWuseC7xDflU0L3QfxnrfmGLBIgPsaEOpwZb6HiECt3TP
rZY+XdSkH4lY6omSSWNTV2Lw8EONRTiCKVwTP1lZJpXFi5iCRQI1fX9c8gM7hiRG1XLlnx7B4GwUy0XGqJX4WwfvdHz69VGv9dDKMywNO2nCeGlVO/DCgmv9+0YTEOIT
KjSSNhGh9eaWp2daon/nCcBOcKRSNrPco1YF5pwPwV/nni2uiPG03BOTqTDCBQotCr375Xs3tNp5P3JQuDF/euNRZ3wnmZBSZmicGpVWuYRTpuA7aHOlUzvSIMDFGxtb
xSlXj8SQxMV0eMt5mwkUCLLhoGOLpatml9mCgyzNYSP1l1HW17IJewglN7OmaEzMN/rDrh5KrBCleDhISTJGrUlvTRegigbhy3a32fHRKvZWfOtbGW2RMP7K9pHDhFTT
w04ZNB0m27sv0riZEJG8aeu8ga6b6wT/6uJE/xqcaiXL78oFxG/Lp76qf+XkryUKQw3g9I9xQ3lRpTdaraWrWuseC7xDflU0L3QfxnrfmGLwY0ewB+Px/2tDbaLFcrCX
BBGg2U7Y8NtatL1SYWnXPcj+T5P8di6XieeA1YJl3fqOEfMyYXt5HPmQF3upyAS2GjiCMGxE+Jhb43u6l6y29SSNhsneWrjn6ocLnmeTYp8GIsyw4PizIlx9I3dyHY9i
iqxmHsql+VujH4ayoWS9r20dJMul6zgeHMxKJ7hLkYr7DdNTBouIDyd+0h5pIKvKgWe1eISIbGlSTF7anQaFHHEwwsNttwTmcczwBsuVGnEo5TwLj9r7KUxOXC4JBh77
htI/Vu8MJaYwqhb4WZAsFPYkYrONHeYqsSXreAo+AwO7bs+NlNQF5CvKlWMj+5YdmPParPwu3NSDIxzC4/LKNJoGCa5kSQBKDk7N9B5yBeYEz7OH7NQB8S0bGD5jOdV7
4qJHZaPNRMG+vI8+0H8+UkqL6eb9UPyHPHho0lUh8eSzT9htMgDXbFlWg6dmdkez3A/PxgQYWgYJCytdn1VqUUSuqtFaC4ssy+ITOZpmGMe/l7nlr/mlcamM+8eW2AUe
bb0ZvhE+fOZNNdn4Dk8m+97YN+iWSI0zfA+1UPUf1bJVIefREUutdM++DyhXD0IqLnHKUJK6/DIjgxareYH6z3LTnsWnLgQyGIRydBAaET3fHLQVfYgDiZrJ8boiCCTm
wvKXMgFLcRjXCkEKHfvAWguKWsEvFS+Kl9FGqO8RH6+8gCZW2ghDXdsYo4PGkYs6JWqbhbiJQgB/qil0YMty1P6Mx4JAqrWlhp+JUluLrYCsOBxp7Ockz5a1S2udZx3c
NJHWizosdrRLmHs4SjjTbVbcyDo3EnEqW6y0FlP/434oVHIKMbS+apsVZ6zCe/umSzWLLq88EuSCMnNbkzjOcQuKWsEvFS+Kl9FGqO8RH6+8gCZW2ghDXdsYo4PGkYs6
uZpxLfB+jjyNK1+GhIsi+5oGCa5kSQBKDk7N9B5yBeasOBxp7Ockz5a1S2udZx3cNJHWizosdrRLmHs4SjjTbStm6ffiH7+I4An+57zMTzY21edd5XN/3hBGKeSz/jQR
BAK8jtiyGTjKD0S8xdnAO1MGaha5nLTIlr6IZcRBn0UrueUQm6bSLu1lTx17surfwdBTD/s6LMpMggtF1i1tuDR/oh53SoJMAsUaIXmxsb/Ujtq8y2CvINBje8Yenfas
spgc1EbAyNk0QfeJEmgDVxWdne0500DZrSfKeQkY3oi6/3es07fnC+88jlV6iOzQRK6q0VoLiyzL4hM5mmYYx7+XueWv+aVxqYz7x5bYBR5tMMuN226dJ/btcAQiufha
71BFeVsA7K2EsdtazfFyjWLw8EONRTiCKVwTP1lZJpVse+BqCcjvVxI5s++8i7jh1ObC4F12xIniJ/vPBf1lZuI4tWUfFltSHSTAAl2qG+DR5ShRIl94UvBsC1M5FJnJ
/pSHMoFnljdB86Srl3rzZQLHCtasGnFDY8vYmqi+5GjFiupUpkrgBtPqTrrf311BwnhpVTvwwoJr/ftGExDiEyo0kjYRofXmlqdnWqJ/5wk+t3Gadz6l4NKBsDP4mNCk
OphwATLtaA5C0EoIoK1V9LIFNhX4fE0iGrgbx+h9IiWAFRcKFBbiOT1X/jSJQtiNSW9NF6CKBuHLdrfZ8dEq9s4RYzmqCKf1d4pxbpXdJypx4JXyMEx4hPm7X5qyRayJ
PWSC7M8w31wGGEaPXd72mDR/oh53SoJMAsUaIXmxsb/Ujtq8y2CvINBje8YenfasoNRUUUMu/N806tC+flOd90HTrZOEAYm0bNasVZfEXecKDLQ0qQCNovUuexI/JyB5
KjSSNhGh9eaWp2daon/nCT63cZp3PqXg0oGwM/iY0KQ6mHABMu1oDkLQSgigrVX0G+0XrBhlHe9Tz6855GfcGVA6uSfJWcRYAvcWI279ogCL/s/x7sRLJ8vKulhunbhi
cV4ORQ37S3MgpIOzFn5AHDb8odXMguYgQN4T9epZpjqtlj5d1KQfiVjqiZJJY1NXYvDwQ41FOIIpXBM/WVkmlWx74GoJyO9XEjmz77yLuOG32jVw8+q6jSyf0GXvz2a5
oP2nlh5TEcxZwvL/gIdisOTEx8AjzXJ7P2jEV4w2xN7nIgz052WWswq9py7tYm8LFeuxK8N0q0pTwYkc1DpfLv6qAXEbAokprPsGEqbJOkC0UQPWTiromLGvyNQ706vd
wMMBAw0duLRDbA9vyI+EOYv+z/HuxEsny8q6WG6duGJxXg5FDftLcyCkg7MWfkAcIqeLZk7r7eua92aXU5JOxuOBSNMNsqumGAVuORtuu/ndj57hhMwOPJmJyv4km1Yf
i/7P8e7ESyfLyrpYbp24YnFeDkUN+0tzIKSDsxZ+QBwip4tmTuvt65r3ZpdTkk7GwdBTD/s6LMpMggtF1i1tuLIjnkSgQgSiQM2MNRMJv3nUjtq8y2CvINBje8Yenfas
oNRUUUMu/N806tC+flOd96xffOcbUXx3rvo5iBH1PWzS1iwqrrujB5umy64I1qqDyijZh8LmwfiKibX/WkCyZNSO2rzLYK8g0GN7xh6d9qyg1FRRQy783zTq0L5+U533
xyLPVIXSAl+68/kSuaRvmqoO8NN6LFd6t/5dovnm6IjKKNmHwubB+IqJtf9aQLJk1I7avMtgryDQY3vGHp32rEkilU31mFZOHca7r6qD0CkK41IaCDDFXJQ+j1FRAEcr
0eUoUSJfeFLwbAtTORSZyf6UhzKBZ5Y3QfOkq5d682V/2688GNmNbT8wwMxmchI7lLmHHUT62vSmMdpZ8F/quWxCVpCpe36M0yt4g84S+LTnIgz052WWswq9py7tYm8L
vfsXqFavtQNAIEuAKJWJhD22akT4UpcL8LMiFAamf+xt2hFLlc8LQ/Ink0BJ0rea5yIM9OdllrMKvacu7WJvC737F6hWr7UDQCBLgCiViYR/owcF84fdzg7I+2k/z36X
yogm0Sa9h4GMq195YwJtiFOm4Dtoc6VTO9IgwMUbG1uw25jugxLWOli9ksKqW5ZuUDuj9BX4uW4QIiYSky8Pvmcd0A65H8IyvBNa+olfzXPKKNmHwubB+IqJtf9aQLJk
1I7avMtgryDQY3vGHp32rEkilU31mFZOHca7r6qD0CkDHwT40nxrwT9mr2MEZT8h5o2GRkz6ceXx5Ax9dmnkxlOm4Dtoc6VTO9IgwMUbG1uw25jugxLWOli9ksKqW5Zu
+slIj1F3sZr7K70olxIuFnZQKrKRyBb9Un6xJrR0waYq/NG/OQFjdXnCdVe4ITZsUwZqFrmctMiWvohlxEGfRcIi+GnCvbDdoef+We4hKWodk30t5AAt1T4iqqufsUWw
mgYJrmRJAEoOTs30HnIF5jiv1LeKrhWbmQx/DmJNsMl3NhFJimsRasEAGHoikDVHyijZh8LmwfiKibX/WkCyZEdQMLzo3NB4UkPb7Hg7we4LLFLaTFxY73WsApJEEiuF
GvH95qDuPxUfKLWztzmT0GTcj1vY2XA04YoKEhh4DPrTERIO12COYKabGTFtZBCxfuaM3Ayv1T+p9TuF9iY37b2Phv7ZbKtCltOima4yArquouzwdWtjCt9owoXxE5Q1
coXQKxQzv1NURAi9QM4nM0q2qUlKZVFpnMWiTRCiuFuut0sncEmy1OhuK5vpOZi4pElxVHX5OZBoKwXu7Mfb0huvFwZ7uF76p65+MYtmN4h+5ozcDK/VP6n1O4X2Jjft
+XCwEZo6D3/Cl4TkimEwc1A6uSfJWcRYAvcWI279ogA9CcasTAb/rTo2IKGB4WPBMWJn/U374nmauItfuJWgXhSIcpGCatFyUYstJew1q/XVuHZqIZdnVDqf8SmLU2Nq
Jz1MjxVV/HCqTvskm/mtyNvBKMU5H+LNw8FK2KSAkL/nfDefwRynsaDsu10PNKpBuvvcdE1NVPtag2YEeUjIXiOLseFWtLsqSVLnUox13w0t1D8VXXx3FA92dk3wDiOb
k33xY8sj2NCXod1KWQj0AjFqS9OUW7c3eej3Rc65uaXCeGlVO/DCgmv9+0YTEOITqQpJvmd5aNDU6ls3WoyKWXyCAngh+4+rwr10GmYD0ZDkxMfAI81yez9oxFeMNsTe
gNLWKOrT4wpEWz+2QeXg3Xc2EUmKaxFqwQAYeiKQNUfKKNmHwubB+IqJtf9aQLJkDLQuPz9w0cv3DehpPzVC+3EKFurvijIePthr7258jfnjrfreUw2gNJbq1rtDHSGD
UZ8q+yz32SQAWUEBzAqfBiYgCFm1Qpbz+Ovn79WIOYG/m9ncnkZ7Y8sMy891iWCCUaLwr5BdD5vS5yulP3+e00bxtkYKqN5x7+D8WK+9SZ2pod2kODkB9lHFKaHl8uwT
gBUXChQW4jk9V/40iULYjU89PnhFFBuPLMbLPW7kqz1p9x/TVikdNR+F1KSEHESYFbfecuNhQ8VdgysgNNya83Q6V/rKBoOrFanLIoRf4YCLBQsXlg7+6jxSUEou9ylZ
kqJRANrzttwecA03XG0O3wWmsXj2ah0jEAWK/qPR0lVEx7SDuyF0S5IAc1wGiFcJP5hAMT0F/0AAqXSP2eu/Cv7xOOtXmQRpkqPebs1heUve2DfolkiNM3wPtVD1H9Wy
oANV0IAbPZCnkvEsXCxLHQrjUhoIMMVclD6PUVEARyvR5ShRIl94UvBsC1M5FJnJWvsziXuj9xziKLk3Rq80HBBL9mFYvXCJjYl0M6lfezr5Nys2CawAwRi09+EzY6mn
d7KZ2fLHsQwwei2++Glv4tyqZZUlhITuObGJtSkEgWvZz2yLCprevq834y/XcIgO3rdgMwHcs5xHKxXHDvdw0K63SydwSbLU6G4rm+k5mLil6ZhoEWRdCK/yw4YXJMm1
5MTHwCPNcns/aMRXjDbE3pLKQpkDwkcQf8KlG6wH9eph4YAPvw4jNAzwO9MVn5FF4YkYbu3ZBdgTCoGF51Hy7e3tw//Vo9JWn/tzTMv8949SDUB+nYRgFpW+ojyXLg4H
wnhpVTvwwoJr/ftGExDiEzvIR/w5vH2w2WW/xJVclwuAS4Bxbh2FZhj5WZV2bRJNZu57g17tbF8FcoohXgWVjuCsCD3UlWynLeS4fDBjEsbkaDRMoeUog81+PEF/MFkl
+T6u0B2WU+6gZkSPUOohuLghTLUKOfG0Mwap6LAuGEHHVJusz4AsDRaPSvedTc6T7e3D/9Wj0laf+3NMy/z3j/SaiUDylCl/hCGI32kPuQ26/3es07fnC+88jlV6iOzQ
VjYYvNlhPzr0PoHUOztllGyoExnkgn26/Crp+Tkkn5PYG8632hZu9Uoa15VJKNy/hEIQGK0yWnssnyQyK3jkSt4L4k+UZvvuAPmv7FtuC5fTbQd7Cx8I1r35LA9GUGLY
SWMkiVpavql1mSUfD8Km9EAPjcsG5V+CsAumu/zdHmkCrKWwkulLNin5DOn9ebhX5G+yzcwjohfR4AJqeF5Uz23aEUuVzwtD8ieTQEnSt5pV2aDBLZgTs/r5rAXOydpv
HLWEOhfIJLXk72VRryY1GmTFUPwtPqLVJ5eRwjIxq+PBkN21+2Qq+l3BENbCL8ARBBrFAGOYrl4uarK+eCfXghohCr7VgRWsxxwAmB9PQ1pC2SZ8RS0ftOftsC5mfZf7
yPVahDH1kBucyxt63pxYJiGoB5ZjA39baL/KRjJpVzBEfQsOGD0C9UW3YUF06A7CbEJWkKl7fozTK3iDzhL4tFXZoMEtmBOz+vmsBc7J2m9hNbq74+M7aE7TrRa+IXUm
LdQ/FV18dxQPdnZN8A4jm8dUm6zPgCwNFo9K951NzpPt7cP/1aPSVp/7c0zL/PePGYimOdVdKh4xKNFx/Wn2Pd7YN+iWSI0zfA+1UPUf1bKf57V5hGbPEjYgFY+1Auvm
Mr0Nc9JW4GB9aNApi3IGi6FulHV7eqFl5FOqhHSX7aWaBgmuZEkASg5OzfQecgXmjQxezLAs8fWMyykcrQSAdyg+vrW9xFhmrvHetGFVZI5BQ6pV3Sxaqx4kt0M3P2tw
mgYJrmRJAEoOTs30HnIF5o0MXsywLPH1jMspHK0EgHcoPr61vcRYZq7x3rRhVWSOUd9i7ZhK4KlxCYU+yf6lFeCjrbOm6qMfi3YL8s7iuMyNDF7MsCzx9YzLKRytBIB3
KD6+tb3EWGau8d60YVVkjvd0/jV3G40uCpk175qyaLWEQhAYrTJaeyyfJDIreORK3gviT5Rm++4A+a/sW24Ll9chdOHU/fp+Zqxg54D48QTB0FMP+zosykyCC0XWLW24
rqLs8HVrYwrfaMKF8ROUNW/bD9Of8txvgB7S2FMwos8L2PiTeY0aKnmiCqHbAHg8VahJUgliMRUyZZH4sOfpc5IdCIJ0ylSHFRJawVFwL0sEGsUAY5iuXi5qsr54J9eC
MuhZkpbRVXqW7/FSVRKEIp/e/J0i3NN0SKQJXyqSPm3HVJusz4AsDRaPSvedTc6T7e3D/9Wj0laf+3NMy/z3jzEJh8C7GSl/RBy/bBcQH6QBH2t54ZS6uGvR3/qKOCLj
SnO8v1O1AXS2sQQAaspt1Bbwv3MrNDdl4t4wD1KcBQp+tXdFKQCVv+PSoJRmeCcYOpeok1I1+qBzUkkSmfKCLEpzvL9TtQF0trEEAGrKbdQW8L9zKzQ3ZeLeMA9SnAUK
beYGJUCi66ZTy/2IxMEUVe92pP+koWQ5dxWSUcIA82T5FLb36BxHbTLyEg4Ez6/Vgjaj9K61Zs/n+tKgzF1TpwTlcMjemi7dwTP5/PhUbcXvdqT/pKFkOXcVklHCAPNk
+RS29+gcR20y8hIOBM+v1YI2o/SutWbP5/rSoMxdU6fcwawlYuhOAgLe0kO14PnhW0mjlicR8+7GPaf/YWtCMMj1WoQx9ZAbnMsbet6cWCYhqAeWYwN/W2i/ykYyaVcw
Vyt9mPVIuxBHISRWhSFQkLeLaJ2f7j7IBdYIP23B/Ks7yEf8Obx9sNllv8SVXJcLgEuAcW4dhWYY+VmVdm0STY1Kp5A4h03aRWEPp8QxPDnCeGlVO/DCgmv9+0YTEOIT
O8hH/Dm8fbDZZb/ElVyXC0xlgASglVBJCFz31xAir4ftyUsOJD3CS85a7SzIsCE7y+/KBcRvy6e+qn/l5K8lCsxPknYEKJaKxCEebFgKOgfec7pqvMCVdgl8YcxLCISB
cQoW6u+KMh4+2GvvbnyN+TvIR/w5vH2w2WW/xJVclwvzg4hTw78DwgNHc/wyxIrVDyZ/ehca+67e2ay3GyhP0SjlPAuP2vspTE5cLgkGHvufMcepmSGw/pQn+nwlxBZO
kAGqLX6cih5u7pIkz98Vo8qIJtEmvYeBjKtfeWMCbYioLwU3xOmcT+RUsimY0qQlwnTmnbZ6PO0DF/awJoSunAQRoNlO2PDbWrS9UmFp1z3hiRhu7dkF2BMKgYXnUfLt
yQURs9dieInI65AkphswgEMj9oKWdA8UIw7Bdztg4/njUWd8J5mQUmZonBqVVrmEqC8FN8TpnE/kVLIpmNKkJeCbcuv5QOyOjnSe2Jl4HBMJZLii03xa0EHdK67y6+IC
N/rDrh5KrBCleDhISTJGrWhmExIgztZA2Y3zQpttD4Mip4tmTuvt65r3ZpdTkk7G7Hq4rwJaUqBPtDzIid9GeMvvygXEb8unvqp/5eSvJQrMT5J2BCiWisQhHmxYCjoH
ScWV3XEEuHVocB/RfZmm7GHhgA+/DiM0DPA70xWfkUUVt95y42FDxV2DKyA03JrzyRHdj65vVSLIbvB/fEiWmQrjUhoIMMVclD6PUVEARyvR5ShRIl94UvBsC1M5FJnJ
RsosYufysGc6pDn5EQkm0LyBOiSEd8L5gxr7ugDu7pXTERIO12COYKabGTFtZBCxTAA290DVPuqfHhQ9515tr7ATYqkO2wikkUNA5yTHtNJEx7SDuyF0S5IAc1wGiFcJ
f7KKOJEKqFjITPL2FMfT0TkKD9jCtyk2GTJBqV9Lhl/iHj0rTxoZ6bRub8ATr+vm9vuus5H+VJNn+frGjkcW7qmtAxvBqmFlO0ATy8GPLY5BQ6pV3Sxaqx4kt0M3P2tw
mgYJrmRJAEoOTs30HnIF5ndf3W4tS9jkUXMB141eH4TSd/apBaBrxsxREpUIgQveoSAe+ozQjYVkIfKt0wh4xa63SydwSbLU6G4rm+k5mLivAeVor55mopJjpJWBDLdX
iCOvqWRi+6mWyEsD5GTBndu4yTnHIQM/Be45Cw5HXypGyixi5/KwZzqkOfkRCSbQdJL9T8BXG3Qh+alHQnlrWClZK4Jfph0C6WJsD4NGaZD2+66zkf5Uk2f5+saORxbu
eJdHAefwGW5tqAWDuCR95qo5wc1NRvJx6R1eYWvkB4HKKNmHwubB+IqJtf9aQLJkYREUkbT0pc0v4Fp8HdCj0OGdkjlIuQvKjIu+stmKKZ3KiCbRJr2HgYyrX3ljAm2I
72x90kb2qvC0Qvv0Q26ldfKG73kgIEA+CuYJFUR5kdOtlj5d1KQfiVjqiZJJY1NXRvG2Rgqo3nHv4PxYr71Jneygv8WFy88XcQsMI0jClWxp9x/TVikdNR+F1KSEHESY
FbfecuNhQ8VdgysgNNya85HRndBTVl4YvJIcHDKrGHnr7YGHIrBw79ZVXMMfc9jPaw0O3gjOdZpyp23w0qXyIy1ZJnYR83s15d4MFW6GocmYGDYQudJXegft0Wpnj1Sf
X53apfJV3s12ljNgEiLTxfnuzyvnERQqz/fAmbwDVDSeyx6GURWOQj29jrgXBsop/ozHgkCqtaWGn4lSW4utgPnuzyvnERQqz/fAmbwDVDRR1wULm8FKSPqWqyVAu7m/
DaoT8A/UVctujU264+XwRQ1t4q8u+fJk5s/Hl+9AWoht81yZKbj096jwMruROtzulkfiVouvsklfgOyR/fbyHmJfBKqk058fiWPwO4bGZBDnX8V9sC71e1x5XXeDPIv9
KFRyCjG0vmqbFWeswnv7pvb7rrOR/lSTZ/n6xo5HFu4qyvZwwSf24VETvt9r31gjMWJn/U374nmauItfuJWgXhSIcpGCatFyUYstJew1q/UWnLHnwGeMyHACf2qBVSmn
NYatGyygIHWdVxG165384a6i7PB1a2MK32jChfETlDWc4narxzYqqc7mkZCId4MafmdRDF2vkXSPGhz6FkNRGuwxYcfm5JQJ1VLe5bXzen1VtUUsrchJD78lvRUWXLQu
AeGLMO44JGwbze1ZynvNEubbKrA+OU0N2fHXzFVl55b57s8r5xEUKs/3wJm8A1Q0/dX+c4JcFwWKuSjZlN/lr+TEx8AjzXJ7P2jEV4w2xN7UJy66FSKqpKkQn5j2fqnS
RtuYvBCGgshDpd0HBeDcYN7YN+iWSI0zfA+1UPUf1bJiXwSqpNOfH4lj8DuGxmQQGONVpWLEijtUiXriAXDnMuP9uRzUEnHTeJuWizEiQUzrsK1wupmEpoCynz/bdPSg
QZfL9JOtJkgBKKVxkk+zAkTxqpWR5iankpnBHUHeBctRDdFxVUu6jx/wD8MnQU6xYl8EqqTTnx+JY/A7hsZkEOBlDqC5lh0yACy961lqLTgXCQvYy1mKyp3j/jM2NBCM
XDNImikGHGfIQQ+VyeVpYw2AUbE+EFMeiYElkfqezYjy+bauMXc5BGVMQnV2NUIIuvvcdE1NVPtag2YEeUjIXqeudDrtgtZCJYXNcJE9ttbsVbSVnL6gZvxGRwOUgiLV
q3J1SjMH1k4FLkVcmJSM3RSIcpGCatFyUYstJew1q/XsTDX/0ttuajkEoASeyCGHMqHQXL7OQWxIJzEW38u38ubbKrA+OU0N2fHXzFVl55b57s8r5xEUKs/3wJm8A1Q0
to/MLlw4xzCGUJBuQnVOhyhUcgoxtL5qmxVnrMJ7+6b2+66zkf5Uk2f5+saORxbuBCMPvE83AtaALsU2vNCP/JvWzKxuUVOjZIGsohMY6E5PfGW81BJ69qcC0AKxmK6p
JpptyE0+Uq4unlcNdOw3TTHRwIkaod3gwgFJaG/gPxQKDLQ0qQCNovUuexI/JyB5a6h8cmvKjiIr9+uHvW6/VIEdwQGffOhbRac0JMCZmb1V05QvIgmRHf2aHiEWXtPO
3Y+e4YTMDjyZicr+JJtWH9MRz8Y5Qm5E8uVDfiEPmx5qNR3vGk5u12dbOD5sbYR8kH+R5iaAROlsVfKBgS07ag1t4q8u+fJk5s/Hl+9AWoj2SRMqS4uvynXZBRiqGJdN
YeGAD78OIzQM8DvTFZ+RRRW33nLjYUPFXYMrIDTcmvMxWAsS07mFgl54MSZY/5eNWrCg56sN01Y7cWMDY8p799MREg7XYI5gppsZMW1kELHOKiJaDXqYCm6qPeSA53BS
PCW4/NuATcSV/cdCEJZcJKtydUozB9ZOBS5FXJiUjN0UiHKRgmrRclGLLSXsNav13mqf1mKaEIjwnLFVsGZqBclTRT5en8ca6fx+3IPztibkxMfAI81yez9oxFeMNsTe
1CcuuhUiqqSpEJ+Y9n6p0p2+dzoGYEwMDXQG0PSsSgMG/sr9R/uLe2WcGA6D2ao5yogm0Sa9h4GMq195YwJtiGJfBKqk058fiWPwO4bGZBCseWBPJhGEl15zvta7fjzV
jfh4Ya/9Fnkr/yVkRU9wldMgR8R+6jwHBgXUaTBBMsNG8bZGCqjece/g/FivvUmdju9a/ozOKvEV1DVUpcONorh2xNbB/9Xo3/bgtUcWlguAGHT7EEjSmupE4ZxsNeI8
X53apfJV3s12ljNgEiLTxfnuzyvnERQqz/fAmbwDVDQGLo611ZYaraZjIMtY1epAnEUt4UJjmgYdYVoHUzMRHjbV513lc3/eEEYp5LP+NBE8UETOf2CDlUB9xpBtxMPv
CFAAbDHf7/zBuwSZ1RYjBr8EpwjOLNE6Ae09iMYIQ63p+r/qtw4Lcs40BTF7nYqT3A/PxgQYWgYJCytdn1VqUc4qIloNepgKbqo95IDncFIWf1j7OYN0AOR3Gpj6P4ys
SRyKcA0MDx7CyPd+TOgonTQZV9E9BW9djVSs3NzV4IqSHQiCdMpUhxUSWsFRcC9LQZfL9JOtJkgBKKVxkk+zAkah7Uq8pNH2ZB9YfhxaP0COVeVEOLT/igVMf7IU8+7U
vY+G/tlsq0KW06KZrjICulwzSJopBhxnyEEPlcnlaWMNgFGxPhBTHomBJZH6ns2I5NjecheY3JPsioHKK53E61m1uIlIdH8cp+1f3U3SKWx3nkTVDdP/BK37bzzMZQsK
yijZh8LmwfiKibX/WkCyZB86uSOiJatsvskisszauJzZOh7+QSJTDSdJJELDRp1qFeCVMxCQk/puuMmnIx2dkmn3H9NWKR01H4XUpIQcRJjJ3CP6xjn0ZfLv7pv04GCk
frjw8qipVgsCqoyeWa0GXqVW5tKUtv8WCugypYyBVfuAXDaRR9dUOBQUyaCK/+3lq3J1SjMH1k4FLkVcmJSM3bVFlk/G1gKOA0XiFGMYEB2H+Qr8TcUehGvK09xqj+SH
linxHmI7H7/VzkpfTqR69LyAJlbaCENd2xijg8aRizpp3lo0a1J0hEzy2LVT83uoQbV5de0XGq0UmAe1pUQao/AUubkiQyO9B3/cBfUJmOqPW+wpuBD+vbfDYFomlT1U
PfQ1bFYXDIHPzyXnnaGhC4hGMEqOThYPO+sQ89+UNmPcD8/GBBhaBgkLK12fVWpRONBoNjc1vZS/sPIlWzJeyJvRge5FXjqgYeioumq4dFsJBYOiX5QBLQcd3I9rFrEO
LW53280uqMkncBzWtNEdFNMREg7XYI5gppsZMW1kELE40Gg2NzW9lL+w8iVbMl7Im9GB7kVeOqBh6Ki6arh0WwkFg6JflAEtBx3cj2sWsQ480K2AQq0gYNNdg0lPM6RF
WDJ+cyBSpbvClTO6IEId5V1R8yqDM078dDcdDR4Hs4jAXGeWmG8DVA5m6dL1HzeQJVKa5rWhGmJUyc4UEEuVCBRGEWETBTb6n3Fgj4NWf7Gtlj5d1KQfiVjqiZJJY1NX
RvG2Rgqo3nHv4PxYr71JnepPwD3VVOcZ3V+uvPmsEw1o/HsIKoPXZSUD8jz178XWmgYJrmRJAEoOTs30HnIF5vnuzyvnERQqz/fAmbwDVDSEf4gMGLmDPttk485/mk4G
0yBHxH7qPAcGBdRpMEEyw0bxtkYKqN5x7+D8WK+9SZ3qT8A91VTnGd1frrz5rBMNLqL1jKdWJoyZtvvfIS5mV4sFCxeWDv7qPFJQSi73KVliXwSqpNOfH4lj8DuGxmQQ
T7evWHYuQK9h5P9uTYcYI4hGMEqOThYPO+sQ89+UNmPcD8/GBBhaBgkLK12fVWpRONBoNjc1vZS/sPIlWzJeyJvRge5FXjqgYeioumq4dFsJBYOiX5QBLQcd3I9rFrEO
N337KRjze2EboJMJyBijn8HQUw/7OizKTIILRdYtbbhcM0iaKQYcZ8hBD5XJ5WljHzq5I6Ilq2y+ySKyzNq4nNk6Hv5BIlMNJ0kkQsNGnWpH6fT8B7NehcO27g2eRlTF
nx+zWXZeuuyRapO2a9M5B11Lkeh+ItLm1SyTT6R7aDhElQpsluQQnp2QfqYr/SXIfbVlsZeNUeNhhka4bZyKogZ42DrBIsl3LL0fj+HZIEHDThk0HSbbuy/SuJkQkbxp
i2uThsmN+MVFugDu9SUNItMREg7XYI5gppsZMW1kELHOKiJaDXqYCm6qPeSA53BS4M03FsFhKDwQxjeCQagMBjlrf2hXCVN1zEJbu2INdUzxFUEoeMepFRr+Hj57zFHI
w4PEHMFpSPTDbPmrmYnYxE8HrEAk/WV5hq3Inon/VDFVTFcJNWYysVpHtG7kevqGCzjWlOPtEuGsP6wjDRQhqy86okyJ61W73cURf392ZC0PJn96Fxr7rt7ZrLcbKE/R
KOU8C4/a+ylMTlwuCQYe+4V3WapRMZ7CVulcsAo1RWsGWjDmCth0b+c5ZUsKEjrzM8Q5b2XXZJxMK3JhWqvBChW33nLjYUPFXYMrIDTcmvPL8+k7ItaYXpDgPBzZNm/N
ZtDVoARsGkRFFKQiWZYpDEq2qUlKZVFpnMWiTRCiuFuut0sncEmy1OhuK5vpOZi4xvcfR1NME5qBjhkrMUapm8hCHPCheslXMUMukcrCvmfcD8/GBBhaBgkLK12fVWpR
ERUGIDzjAGNHZR4Gh8drqkPgflzxiqkg5DdXR5DFwfOtlj5d1KQfiVjqiZJJY1NXRvG2Rgqo3nHv4PxYr71JnV6Nk/hQYukpbOnpHGUAvGU0GVfRPQVvXY1UrNzc1eCK
toJVJtxYkSjW84nDmMO2q7NQjTb/UtPrrVlmLA2Fa/I32AV6NMeXU1ycFUepEu9rQE095xHecGbrNUtbeCSupVw9wH388snso/68fZZaQozHjTTItU+a52dxr3NhbBK5
42OMCSRezWqBo5lmVi37cpDdT2rcUC5+gEQ/BhhH+/U8UETOf2CDlUB9xpBtxMPvBQH8CgNjGacxcgAAInhcz7SJaiF5rTYZAtyACyqVLHhQfyEV9tNF70eDjybb/lfB
9vuus5H+VJNn+frGjkcW7k/Txe0kp2RrQrtoPA1gcQGnTRtrSO38MSIrkrYR7rEvgBUXChQW4jk9V/40iULYjaeudDrtgtZCJYXNcJE9ttb8gSZiHLwUSmvFGO1ad7Ic
sgU2Ffh8TSIauBvH6H0iJYAVFwoUFuI5PVf+NIlC2I2nrnQ67YLWQiWFzXCRPbbW/IEmYhy8FEprxRjtWneyHGbue4Ne7WxfBXKKIV4FlY6x7gZjI31yRgKoITqxgM9j
p650Ou2C1kIlhc1wkT221vyBJmIcvBRKa8UY7Vp3shx9b6iC+mpfU377ZTivyM1P43CWhqmHb45TqHfbJtTaCHj3+iJuIoPVjo8xV5jkhqdvg9DM2h9nUjiJdkNT+Wes
aQebXPadgePQoBXPOhMTTJgx1nI7UI251csIJ+QEaTrcD8/GBBhaBgkLK12fVWpRzioiWg16mApuqj3kgOdwUjjdz1iPZrLPKTuvu1+YYJ0+jNR4rzoIRBhZNkLUBZyE
fqtjCkZyvgTZTF2HSZe8xlwzSJopBhxnyEEPlcnlaWN4PLx/OsERaBadd4HFwDG1tpgnM3ZSMLTvNIzSpRxxsKdNG2tI7fwxIiuSthHusS+AFRcKFBbiOT1X/jSJQtiN
p650Ou2C1kIlhc1wkT221rko/RnJgU9LSHXVdW+wNG7tyUsOJD3CS85a7SzIsCE7y+/KBcRvy6e+qn/l5K8lCi1ZJnYR83s15d4MFW6GocnO/+1kjc2jdmj7CzLi+3Yn
ykpcuO+kuOTpVU/Mw09qmowhdr8MHw5OgArISqYcq1W1wz763vulT3mf0ItXqIltITftZNRlXFQkEde4wrxDwlB/IRX200XvR4OPJtv+V8H2+66zkf5Uk2f5+saORxbu
kleFRDTONH9rEnlyIPluoP3KXbzzWgjRzrCGczMJsyC6+9x0TU1U+1qDZgR5SMhep650Ou2C1kIlhc1wkT221hiynBURXuKhWBWMziqkT+rYG8632hZu9Uoa15VJKNy/
hEIQGK0yWnssnyQyK3jkSlW1RSytyEkPvyW9FRZctC4yl25WTw5UKkKPGn/CWRIWfxcLnQylypxZnRLmA93hsBSIcpGCatFyUYstJew1q/XEH432QlsiA6rZ7tAns5TC
nmSHeCltF1Ci6ebiDRxK4St4yzJRwMwbtPp+vPYF5BFrqHxya8qOIiv364e9br9U5yBClhG4PliWU/t4d2tGFZ/ziYX8Kt6Sh8muutkQJp3NLBK42KSKL0/e7GM2D/ml
zioiWg16mApuqj3kgOdwUmIskL9N2liw4AnrfbwfW8SjZ+4MzfLK/DbXPiSYSM1g7DFhx+bklAnVUt7ltfN6fVW1RSytyEkPvyW9FRZctC4v74xddJxSdfXCYIWrF7G9
COPwgfSsfykNqo5Xvbu6Gq6i7PB1a2MK32jChfETlDWc4narxzYqqc7mkZCId4MasLabjVIp+H0v7JCZ/37Mp4EhFAYoSae30I2gFsc9QvL2+66zkf5Uk2f5+saORxbu
kleFRDTONH9rEnlyIPluoNKy8ZRQNIcB48iHejuvksjcD8/GBBhaBgkLK12fVWpRzioiWg16mApuqj3kgOdwUmIskL9N2liw4AnrfbwfW8S0gRNIYYMdaYcw2QxG4em4
YW8JtUeNvgDmhO5YlfwCOreLaJ2f7j7IBdYIP23B/KtrqHxya8qOIiv364e9br9U5yBClhG4PliWU/t4d2tGFXAZW05U5pezozpXcrtP/9hIHMTesNBbH7AqcbEFvHm4
9IW6ChhuYK+SxyH17J1e0LeLaJ2f7j7IBdYIP23B/KtrqHxya8qOIiv364e9br9U5yBClhG4PliWU/t4d2tGFWSjn8WoJ/T+gAjKDshmEus1KKURV5Q8G/uNA14+QnH+
5bUvXUeL+xGlzwcXJnuQhGsNDt4IznWacqdt8NKl8iMtWSZ2EfN7NeXeDBVuhqHJKD6+tb3EWGau8d60YVVkjgzNMsroEcRySSFaHCP+4DVPQtFoGWwx7XPB+1yMcZVc
jJK/PDrPOSgy47mc0tAey3WmMcfHyfbubhvKXa3w+gjTERIO12COYKabGTFtZBCxzioiWg16mApuqj3kgOdwUmIskL9N2liw4AnrfbwfW8TNhXFFCZlL7XX20HLwJGG7
vJYWntQdS+GLDSk4CASek5uMMo3/ykFFcJy/O+hthnhhbwm1R42+AOaE7liV/AI6p69i7qjPkiM7wd8xO8b+3muofHJryo4iK/frh71uv1TnIEKWEbg+WJZT+3h3a0YV
YY8oo6Tmbvg/IZFVRiilvFfks5shxHaoZiO5sBViDUgIbnHQLLqmqPhi0Pdlj15XUPOA1zFeeG1AaF+9jls+2+kQlGAn5DEw5tLLOuDa+/iSHQiCdMpUhxUSWsFRcC9L
bmn9+YaqLl/3K4RP/WTkqdchdOHU/fp+Zqxg54D48QTQDPHPcqufnI6A6SFKBuzGVwsEW5zi8QLpozuuJgWl6xASaD/Op+/rMe3UbKzIhbu1TT6DJG23F8RbpjjXQYXR
ugpN6ETPpj4hVLqyDp2LJaeudDrtgtZCJYXNcJE9ttYYspwVEV7ioVgVjM4qpE/qz6V4OmdH7lpZ+Lz2lQhHXLyWFp7UHUvhiw0pOAgEnpObjDKN/8pBRXCcvzvobYZ4
YW8JtUeNvgDmhO5YlfwCOka6BDNp387rS3IzNKsmJYBrqHxya8qOIiv364e9br9U5yBClhG4PliWU/t4d2tGFSXJNuHLUqDT2PnuMz5c/8pIHMTesNBbH7AqcbEFvHm4
ET32frxKSSoWfOoN4KNL34mZBrOwHf0y603dAx7Y0rjDkHnnN5oK7j3+mgKZG4QeaNjASzpDNyVtWCbpPyGfwpzidqvHNiqpzuaRkIh3gxqukod4N5FNqjvegS2y3isF
5GsGSZg1/WTNHNbrpTMnjFcLBFuc4vEC6aM7riYFpesQEmg/zqfv6zHt1GysyIW7tU0+gyRttxfEW6Y410GF0br73HRNTVT7WoNmBHlIyF6nrnQ67YLWQiWFzXCRPbbW
GLKcFRFe4qFYFYzOKqRP6n8S+AWHFsSUjWhasDLVplHEtFr02dt+u4vIHvXLfnrYCpIZYwQfDRG+3q4+mYAQqKjiEI2jQGCLbjJhc5kZ/0ciGP8sbF0njmT7/2yI8rkq
9vuus5H+VJNn+frGjkcW7pJXhUQ0zjR/axJ5ciD5bqDnplhXdBW5QPULOdN3Zb+hmiMg7hcjhTpvQJqU2j4Hs4P4dqp2+7qizJp1T1iV/hp++rOM5P/fZ5KRvJNaEtD0
rYpuGvPK9yTRCcxoqu5lgJN98WPLI9jQl6HdSlkI9AK1wz763vulT3mf0ItXqIltLMfNmgnytZxPHiKGyziHDsXPDkT0LFCeSSTzVPci6Mcs+F7mu17uP/jRgWsyx7FQ
+g95P7urU9dWfniP+g400kqZxSgmLt/I2IGp1XcjXPqaBgmuZEkASg5OzfQecgXm+e7PK+cRFCrP98CZvANUNN5b6tDFtNM/4Gd9G2x59cq5XBLSXxgX8HIzaKLFlda1
vJYWntQdS+GLDSk4CASekz7ga+gs4rQX1rZA2lC9ZXyaBgmuZEkASg5OzfQecgXm+e7PK+cRFCrP98CZvANUNNAKNE3ttfGNvXheQw5llhzyw83hJU9bEvbAexr0pSkE
afcf01YpHTUfhdSkhBxEmBW33nLjYUPFXYMrIDTcmvPL8+k7ItaYXpDgPBzZNm/NjzAX/om64ll8LYWUeSB/HLJ3KT+gzh9BvIv+8LC5IMFxChbq74oyHj7Ya+9ufI35
a6h8cmvKjiIr9+uHvW6/VBJk4FwGxXhLdm+DlWOd3U61cCuYy07pmUyAD+5c350TKFUNu9LuhPZqlbgV1Z61ThzvqMthay8m/8q5U4YIdl4a8f3moO4/FR8otbO3OZPQ
DRJn7QKQENWeVPHYAXBM+0KVWlyka/nqcCTbXen2pcPSefamXW7VZEJAgC45f8mcKkHTYLZ3eFVgR6Fcq8b8rPTqStWu3egU1M+KoJL2NVpvg9DM2h9nUjiJdkNT+Wes
gEGBK7tqZwsDqep6TCNDF5SXX67u5XthD8AJQL4/BwuqDvDTeixXerf+XaL55uiIITvOaUXpn5wp/GySvq+pzNFUwEv/cRk6CN9tEz9jtSlHbE8R0jHvFGkRAPbPyPGB
2nxSsvPvV3xnK58zc4otq5S5hx1E+tr0pjHaWfBf6rnoLrmcMTWgL0cmb1rtUAU4EUiDA6G4NtARy8Hj0JVJQ08VkE5SNQvAY1Mih8waGeI8w0agJUN/6PzQcnO6Rsj6
llRfZj/971AEh26BM7MqP0THtIO7IXRLkgBzXAaIVwnf/AhDPr28zG7PDFs/FGcjko6r2p24EFGxD7vAKUjai6x5YTLWaXazU9lvhBIaXNOE5h1nqwZbfc8QzZDh4OM+
NSilEVeUPBv7jQNePkJx/uW1L11Hi/sRpc8HFyZ7kISseWEy1ml2s1PZb4QSGlzTJI2Gyd5auOfqhwueZ5Nin53H8mDXduXrnqyEOSxv0u5j+4gqUBEw7adqR4d8Nhp7
NSilEVeUPBv7jQNePkJx/uW1L11Hi/sRpc8HFyZ7kIRtqofDnac/tjpLzwwkzbE5IqeLZk7r7eua92aXU5JOxl4EXcjCUVETucR0L2XfWTJQZiUf/B1iXF4oNGkYzJN5
mCRSRBsIE+Js0S2ABNZ/yhjzTbbtcRNNFKamzAJ8kRTcqmWVJYSE7jmxibUpBIFrEdLwbeuTdWjTa7jim1RvG4gLXkNKejMLtMzt4Wi6+5cBrqed4qgeI3OCJUtgTELW
bPO8vx950MQrn9D7dzPKSOqk6H95cxp8MXIpC8g7SYFEx7SDuyF0S5IAc1wGiFcJ3/wIQz69vMxuzwxbPxRnI+KXYIFS891oaWKxDIa4LZkOdpRkugaJvOfv2565/h8r
NuHd0tMr+tzC6Bz5q9URR5YZPbxnBIPE/y6kLSq26DpRovCvkF0Pm9LnK6U/f57TvZ+pm+RY0Y9lU1IlD+8R8G4rZvjIiM4afhZgB2ecIzpIHMTesNBbH7AqcbEFvHm4
fmuDksyEc+LjUtJJ8ndm8MJ4aVU78MKCa/37RhMQ4hMbw5CQQU5OxlIzfeyHpUPytOjHwQlT9prK98XHltfEJuTEx8AjzXJ7P2jEV4w2xN6TvpQgS+8MME0frzLXZ4LZ
6+2BhyKwcO/WVVzDH3PYz6BSflgouJUWtYKuG30Ulr5UwwY3NatmdqdtGkC+1mZYKFRyCjG0vmqbFWeswnv7ppi+MDJEOd3C8F0tF2+M2dZ0BDsz2wpFO1Dil8tOYw9D
5MTHwCPNcns/aMRXjDbE3pO+lCBL7wwwTR+vMtdngtk4mzWbxzuHhaAEpN5Cr0HK3A/PxgQYWgYJCytdn1VqUckR3Y+ub1UiyG7wf3xIlpkDHwT40nxrwT9mr2MEZT8h
DaoT8A/UVctujU264+XwRQwokXyLKmuwoSV37jr2myAXzlZflgnMM79EduobDZpAbdoRS5XPC0PyJ5NASdK3mpO+lCBL7wwwTR+vMtdngtkdrRa9zPtIcDlGG2/UGlkQ
k0QdHhJOpsBR9VkT3bsKiDDDX6rfRTIjs9ijnhoeKaOv4eEWLVDAICVg00urxbp9UaLwr5BdD5vS5yulP3+e09Bb/gMGJok9Ay3cwJbYkuyQ9EJIPpxDqBIFB9hlq2Mo
UaLwr5BdD5vS5yulP3+e09Bb/gMGJok9Ay3cwJbYkuzDw3m14bxdFgEQ5cyrGRikXaPqzI2V5ifK7f8NU35SOcqIJtEmvYeBjKtfeWMCbYi4eVuigUYcLzco9OsS0W1+
WRFn7ssBCtFJodEbG+0ousJ4aVU78MKCa/37RhMQ4hMhbk29D478B5pFNt0aSBNDuxzKF4wYF/b3v7WznDlII0d62ZaapOxqmUQSLESSLLAPY8sSqUwff3URBC0NwKRC
WihXsnH/uiQqjX4E7CFoNNyDekyeIyN/9x+N+ecitOoWBAtvpHTa9YyANhLSVJwU/xfrPq3WEj5N3pLA/i+jm9yDekyeIyN/9x+N+ecitOrdJFcvwReiZgZFyk+WA8Gi
7jnuXk6YRVc4bzvYNEW6cyhUcgoxtL5qmxVnrMJ7+6YwIS6gR7C+vDqVC1rXw6qwSFDjdX8TOLPrVAF4oTCTeFvNTIlGMOuwkhmRfOSOtz3EUdutB+iJ3eEuo8FIqI6Q
ZByW+6K4iJwn5FciarTNgSh0ihsCSCcX8KqBgxEOu3XEUdutB+iJ3eEuo8FIqI6QZByW+6K4iJwn5FciarTNgfm/xNV7Ipps9R8fuUpZlu7et2AzAdyznEcrFccO93DQ
CQX5ORxFrcrFVHNCwp/x5DIr0WckXQML9Zk6ehSMffjCz0BiEPTZ+xZbdPRgNavYi8g8XgMVetz37saKphAjidj9mFEnsIrogxSkq84JShAodIobAkgnF/CqgYMRDrt1
xFHbrQfoid3hLqPBSKiOkM5V7pCNszULk3GQkIEZaZxCPI+gjXMSK1xvdhmQoAPqIOG4W1aFTUfJefrZofanFh+/yUqSLUsQLzvg9ldTL2BIUON1fxM4s+tUAXihMJN4
W81MiUYw67CSGZF85I63PcRR260H6Ind4S6jwUiojpDcB4HVb1N3u8JQcQoFDdEWoSh8+JlgzhepTRuZGNxoNFp4yWt1Id0LlEuhiACHe/43KCG5Rq7QG0DlJd7gmmrh
7jnuXk6YRVc4bzvYNEW6cyhUcgoxtL5qmxVnrMJ7+6ZVElRUSuf7GSwU7NJ/gPbMIhbesR/OINzEia76wj2EHr6d9opf5AKai25iWjQ2bSVaeMlrdSHdC5RLoYgAh3v+
YhoPvhA5wdEh1U+YMS2li/8X6z6t1hI+Td6SwP4vo5sUaMPBA1lsVQ12OANLyfZsvXao1P2cAcLQ+DH8qlk/squUGwcXa54CLA5JACBFpgwreMsyUcDMG7T6frz2BeQR
Zmrb+rPs7Nw3EVrY7C1wIQ9jyxKpTB9/dREELQ3ApEJaKFeycf+6JCqNfgTsIWg0Q385kSVAfcyk1nhBRGMg50ySKbn0FWfEtvrkxzaoIqk5a39oVwlTdcxCW7tiDXVM
dIpgDNueOluEswTeNALJsNk3yVl8Kd99Frvu/PAzQ12zEo3WBOEMdIXZ1+4Ek2CmuxzKF4wYF/b3v7WznDlII6Te0+TnGIcVPIcqkLFhlUqh5+Nk/l5icYZwUUyYYUHn
OWt/aFcJU3XMQlu7Yg11TOp6TppMZZELsjOxkAwK7B62RPPdjnNHpJ3MWiMmUDNNNtXnXeVzf94QRinks/40EejWvV5zAnCYwFT2nSbIqzHDw3m14bxdFgEQ5cyrGRik
XaPqzI2V5ifK7f8NU35SOUTHtIO7IXRLkgBzXAaIVwngQvL03L6q9sXmldbtOdZ/LoSEeKgJWnIMlsJbPIcLZTbV513lc3/eEEYp5LP+NBHTNtGeNuUKHKPMKT5OueNj
kPRCSD6cQ6gSBQfYZatjKFGi8K+QXQ+b0ucrpT9/ntMMv8tJvBDYYwigrFeADV2g7VxMRVT38MXHzweO/BeQyJlUCaKpOtu4cBeB1ig1CzTVbIFiPWmzbYogcW+UucXv
sGoRVwU1m/5sVkGIXA+pV6/h4RYtUMAgJWDTS6vFun1RovCvkF0Pm9LnK6U/f57TdqbucSUbn1sDZqIIsp4TytvHmcrc43N4nzZKetCm+eniHj0rTxoZ6bRub8ATr+vm
ny47onHxS3i83SNyGgF8akITTOk6b1Mh6A0hTUofAzjKuXNU2pwmv6LqrVtjsOhQk0QdHhJOpsBR9VkT3bsKiCEvsfzEsaqbEO5iz4WeGFj3hL6gIuleXG0YQ+XRdIjH
4h49K08aGem0bm/AE6/r5jV3toYUjloH2HxSK3cH3iKHArXnnDpQQ62+5Hs+wd7Zt4tonZ/uPsgF1gg/bcH8qzuSByHHx1C9q2vp19yeesToTe9hBAolxnxEVmhPZeQO
e+ZjXMr6WI71uZBbbSbdJFshF7kJQDlKMBcl56jA3MDvCgaoHYihZCzHZVNFBH5C9bcrb2RWxro+3TBailgg3reLaJ2f7j7IBdYIP23B/Kvdb89cmmNrWZ5lPISFB6LT
9iudsG2dCAMxrFMl35ve98qIJtEmvYeBjKtfeWMCbYgwWfcGJqa1Uqs6DSzpymyQvsEMia04GMSi/ypp8l6XIiiuv4Sb2yJvDTVYqhmeBtKeCZnmYzzIodSZyxJptU8K
3AtWH0thgEcLLqWxrOOQzF4mNVSScu7qHq9f4o2T+knKiCbRJr2HgYyrX3ljAm2IGN3ruXPbGFzxk4YHoNL/lbpLbJXKfCC1CafTWghR7pLKiCbRJr2HgYyrX3ljAm2I
cZx1NTcA5FPVYczZ1WdQmO+uChpypypqrL+zthPBtfOUiVNeC+9TFPoxxavzLvxoUY4r6odT1uobKDCn1q0wqfPPXIZHIV6jsjBx4xT6rOMXCQvYy1mKyp3j/jM2NBCM
poHz0bmIJINCoLYSTxpIAVvhVBhPFCsBKwpr9LesuYCtlj5d1KQfiVjqiZJJY1NX0SF56kiHDm4/PmB7mUlb+8VpHOH6IoCNyoJ9FGhkrdpHbE8R0jHvFGkRAPbPyPGB
cDcpZblpBO6x7Q3AQwc0gcIMMSWKbspZUGcXmjYm/9be2DfolkiNM3wPtVD1H9WyZo4fBNbY3dBCxZdysWooCU903/qWB3glMvwgEb7RqagPDjssEpVuHSpP2AAlY/f5
uwOPQ25eSAg3nYe6T2QWQc9mvDIjDoU7ojau+nGehFXq1nm+fF7rd7cgIlvNjXLfs0LuJFF7bZuq6gp0PkAsIqDnvrGFYFHuiqVmmXYrC8syG+GhVkMuf2wU4J3K7Ihy
F9XhIg6/8jOuqWaLS6l7n5p10/jk+IQis4ClCUmMqKb0OjBnBqPxJQfe8pfJ1fT8zr0utT1k2Z8ECR8OCmYv9rmOc/1Ih1KsLB75jq5XqURST1yh09ndfvKYgTIMq+WJ
r99M79Im3PtYEvhrinTStHtRUL2lelZc55mZLAI6V0n/CnAaH1MsgKYIMJ1sBzyakN1PatxQLn6ARD8GGEf79X4P4SgKblRDCNTSKvnYBCuElrw06oPgFCh1+lK3ZuUf
lYVx9A4T8d6a8gbgE4sUO2iMaPVxuyjiyjgiAcTp5Y5Mk7aOs58AkAS7w4D7A0lzF/5dxXb3Bi4hndm4zowyTiJI8WypuHMvD9q2xvR4DozKhutP56KtseqsBQIPMSVz
XTRj139g7yvxfVMItO8P3g8mf3oXGvuu3tmstxsoT9FiUffPP/RpFpYIpIxtX3EsbB17LRMisvxpl8IzgSxptZDdT2rcUC5+gEQ/BhhH+/V/NMxpBCvu243cSjvVWg9X
yfBr5qz7Y0OUuKQDtkAJTcqIJtEmvYeBjKtfeWMCbYi1SJvx2Izk/DOIbS0UNSP2zo17k6edWO+WbLbyfSz/APpcFJJzm9PLAQgzeg70IpCMW6QvUxp/pgn0zrzKQvMP
rZY+XdSkH4lY6omSSWNTV+aU71zFfXofo45ZD+LlHhAiKB/8lqqsow/7J829KwfTGKp73blVz3UUxxPs8JYt5gOo6QMjK/tEfF/H/nOuznrZq+n2onsJCPZjAGb0EMmY
yogm0Sa9h4GMq195YwJtiLuwqqT0nDjvfGzptzrFz4s/QaL+h5gQu7B7aXOWe+sUR2xPEdIx7xRpEQD2z8jxgaQbfo77Im1Pgnxuc6hBSSLeyHgw19VxgLnsmDv+5wtx
KkHTYLZ3eFVgR6Fcq8b8rHWGIWIGQQZqdjL/3osFDPbK2/nnO6BNdw4ME6GofC5CwtuXb2IuyqKqCcW7I7vqcyr5lr5WAt+JAsmNCif5rz3M97StWrZjzAn4pq6oqalJ
bQIBl5Gyn80wkYwHqUHxlBjoxctGMsi2N8+j0FD5yQELyrShRnvTy5qa6oR71dvX6PeWM+ZDu/WXQky1KdC+LJ/4aR9iIhqUzLBjfJYT7e8U9egoVTmB0tPpETx/nGmP
3nZ/ZNweoDeUyZPIwv3dKcJ4aVU78MKCa/37RhMQ4hNsVsusulDl7yBsoL7+wQRiW20fBp1ZreHXUAGQqh8l7JDdT2rcUC5+gEQ/BhhH+/Xyp4Gaz4XiuXOnTqA52ziU
tC6T31gJ9sOwnZVL263bJIxc1mlRW7IeHZ1kM/bNe3MeGmF8ENpoDPMZck3Wp78Wdm8aR3400lRy0X9yOnEsaGYlBPLMMz6Twx9hS6Rt2zEaRS77fb5EyoRo7Faf6zKM
RadI6aAQke0Uy6V1oQrn/U3rFbf+gtNR3MBR8BfflqGf+GkfYiIalMywY3yWE+3vFPXoKFU5gdLT6RE8f5xpjzLPeySFBk1IJMraARxqQYVHbE8R0jHvFGkRAPbPyPGB
pBt+jvsibU+CfG5zqEFJIquG6q7/8OOx2KBWAbbfgWHnXkNVtW0xO65Xi/vivL6QCt8cTP/wLod5NZK/BxHzQmYAOrcfFNRG1LgzLoh87x74WwdejHJrzkldCkg9Pkgq
zQJwZqgzNmUmTaIIYqV1OxT16ChVOYHS0+kRPH+caY8EMaB1mi9rO4vDlku7M35ehqaOARRi7pz9VbxcH5xo45zJCWrI5FVadBTx/FAFj5YDqOkDIyv7RHxfx/5zrs56
WQYOSM5nOpteU4r3mbdH2ZDdT2rcUC5+gEQ/BhhH+/Xyp4Gaz4XiuXOnTqA52ziU4rff6aK2gF1OqpTbmaxyyAXk0LLhtzD8xXNbQ72UV8NEx7SDuyF0S5IAc1wGiFcJ
u7CqpPScOO98bOm3OsXPizomWlv/r0hy0mBV2cZsmWy0F/9PeUVnrMFNCGyILQvSWLw2nThS4rvQnVP/v+JAaYTlv+6lqZRDuGon3/uGUFblyDA2BacDYzwb3aNMxTNd
KkHTYLZ3eFVgR6Fcq8b8rHWGIWIGQQZqdjL/3osFDPb3UfpG7sI3Zur0yKP+bfFYN57XJKa+yJUiKShQrCDVMbscyheMGBf297+1s5w5SCOL0360y0qrLdF3Bb9iRzne
bg1oxkhsBljiASvTje/oS+mcFwGFNnqnVuf5DpT3Q78QfgU61lWBlcu7cC3AOGUNFPXoKFU5gdLT6RE8f5xpj3U+e9StpFjhayEgGT3LMqZp9x/TVikdNR+F1KSEHESY
0Fysf5hhJYG13Klwd66PGmYAOrcfFNRG1LgzLoh87x7xHcH1g5WhunknMRKYPBvbK3jLMlHAzBu0+n689gXkEWxWy6y6UOXvIGygvv7BBGJOaKraJSKZwIl+/cSTgDu2
k8vBzwHoOXZl0GUER3v+ZrF70n3BsRHmaaeIB1odgNW7sKqk9Jw473xs6bc6xc+L07XlGaSQ1iOfsvWTuTpHPnc2EUmKaxFqwQAYeiKQNUceGmF8ENpoDPMZck3Wp78W
dm8aR3400lRy0X9yOnEsaKDidBPmfHgkRVLUXVPXRBYoVHIKMbS+apsVZ6zCe/umpBt+jvsibU+CfG5zqEFJIl6ye5RhH/VmJK618muB3ZsJWWIVJIMZvEkHWloq/ktn
sRfVawYdN/8NRGnvF+x3BYvTfrTLSqst0XcFv2JHOd42ND9CM5kURW5PJC7sbPGuHq0q6oQOizW8Ogox6BYSkir5lr5WAt+JAsmNCif5rz3M97StWrZjzAn4pq6oqalJ
Cmx9cvK9Dm/Dxm2mWzH8gCDhuFtWhU1HyXn62aH2pxatmOt4aeq8RBOHRVXEqram829ez1zl/6SfIOLaOfUCiCVAkXXjFxtzZ+Zp83KbjTs9NvhuYFx3mUy1I0bfoLN8
bFbLrLpQ5e8gbKC+/sEEYk5oqtolIpnAiX79xJOAO7bbUprrOh/pe5vApZTd71feRKryLGHBBi/A9jRApBhHeWrGntEqzz6iFJTXyzRcTMAz3Jgm0AYXxupU2F/X7fMR
3rdgMwHcs5xHKxXHDvdw0A+QcQ98p18sDGsvz24Poc7it9/poraAXU6qlNuZrHLIBfD3gg+nuZ7kErcfhTJW3U728kUeZ7sin9oWLIVFvlOkG36O+yJtT4J8bnOoQUki
XrJ7lGEf9WYkrrXya4Hdm3GbxxQzufpKpzTE3/hCt4kaRS77fb5EyoRo7Faf6zKMRadI6aAQke0Uy6V1oQrn/Y/DgjFLjqr1w0bPqYTxMJbs8zpxvNX1mlF9vvZuZMb3
b2h6CBd8EeQsSs43BReYHvdR+kbuwjdm6vTIo/5t8Vhk/4FXzU0ke87GWwxmjdqmRKtQtfm+6jCvHrfsszAwO62Y63hp6rxEE4dFVcSqtqbzb17PXOX/pJ8g4to59QKI
GxoP9G2auMj6KtDKb7AOuBjoxctGMsi2N8+j0FD5yQELyrShRnvTy5qa6oR71dvXIoefFINhFOmQCKLhuu1J+YJC2K8A+N8Bmwn2fb8A6aUK3xxM//Auh3k1kr8HEfNC
ZgA6tx8U1EbUuDMuiHzvHlBHfRGXzUTf6Iy7SJwUTx5ebJ+lz3gZ4J61woMiX9PpD5BxD3ynXywMay/Pbg+hzuK33+mitoBdTqqU25mscsjI8+BqmX7Mc3OBmSl3KzgU
GKp73blVz3UUxxPs8JYt5gOo6QMjK/tEfF/H/nOuznq+/S+h1E2zrMMOU6+Hrgv4vY+G/tlsq0KW06KZrjICujpyNeLez1D1/xjCx1Vi/912bxpHfjTSVHLRf3I6cSxo
FW9RrL9kJjCVeDob7a4kNjKwnbkZM8pay7kqDDnI4KdvaHoIF3wR5CxKzjcFF5ge91H6Ru7CN2bq9Mij/m3xWBFXDwAgRtc6FRCH0D+mTr10wYg2RvYn/PAGNKEI5xXG
hOW/7qWplEO4aiff+4ZQVoWjVKlFZhEI7dvtWH2vMm7j/bkc1BJx03iblosxIkFMAOge/gzRSQ+NSW+vKD5oFMz3tK1atmPMCfimrqipqUkTuSySp5eweGMVGKmtTMFH
viVLMaQflSZcDFcSiJ1bCjRnRBekJDXEmEZ7MdCWzIt2bxpHfjTSVHLRf3I6cSxoSRiAO8BM/ODFOiRrxPTPRd7YN+iWSI0zfA+1UPUf1bKL0360y0qrLdF3Bb9iRzne
U93+y12Ei36iVH53gFw+tgUrmuDKb2iLYLsO6OmS68pSLc7ePBAS2/aYf9D7fN/dA6jpAyMr+0R8X8f+c67OenpIdGLTTFoPZqVrN37Ra2Tjp0BqVU87LGWDjsZlJF2d
5w2ZhJGrzYh9iEwK8Tl9egvKtKFGe9PLmprqhHvV29fsJUXI0bg9AFlQReiGrQ+EkN1PatxQLn6ARD8GGEf79fKngZrPheK5c6dOoDnbOJTit9/poraAXU6qlNuZrHLI
nLIQ2bBoZtVLVWWGrMsgerscyheMGBf297+1s5w5SCOL0360y0qrLdF3Bb9iRzneU93+y12Ei36iVH53gFw+tv6PrnE5eJy4PyAu332v1aWxe9J9wbER5mmniAdaHYDV
u7CqpPScOO98bOm3OsXPi4cXUh5IttcPDeseZcTyYJoerSrqhA6LNbw6CjHoFhKSKvmWvlYC34kCyY0KJ/mvPcz3tK1atmPMCfimrqipqUkr+lNRSskrXE9+Wp2bDtmP
3rdgMwHcs5xHKxXHDvdw0A+QcQ98p18sDGsvz24Poc7it9/poraAXU6qlNuZrHLI+Zl+5jwL5if/Grt+hhc4XESrULX5vuowrx637LMwMDutmOt4aeq8RBOHRVXEqram
829ez1zl/6SfIOLaOfUCiB0xn7Xizo1lz72UUyjCHe8YqnvduVXPdRTHE+zwli3mA6jpAyMr+0R8X8f+c67Oegu4a9dIRd/4P/tnGKCGEtXj/bkc1BJx03iblosxIkFM
AOge/gzRSQ+NSW+vKD5oFMz3tK1atmPMCfimrqipqUkvLtDw+CwIsq0xWZZRFM/G46dAalVPOyxlg47GZSRdnecNmYSRq82IfYhMCvE5fXoLyrShRnvTy5qa6oR71dvX
TSt4cKHX1HjhQ5PnlwYjqR6tKuqEDos1vDoKMegWEpIq+Za+VgLfiQLJjQon+a89zPe0rVq2Y8wJ+KauqKmpSXGgHCB+Ow6OtzIwWZU4m5Hj/bkc1BJx03iblosxIkFM
KvmWvlYC34kCyY0KJ/mvPcz3tK1atmPMCfimrqipqUk7h1FKwGW7Xpv9aZbiDHpA61HMisGgqrQXJsrgLyGW7UWnSOmgEJHtFMuldaEK5/1FLq8pDQpfNnXVPWj0+Aqb
rsgnB9zSjYueDo1mIF04OblGp9GyyVXUIl39YNIkwOOJNiA9Pvq7uUWFEAMVuGz8sXvSfcGxEeZpp4gHWh2A1Xm5VBrUkBYOum6gYIxmi7VTHRle7p50peXDNripDsuU
4h49K08aGem0bm/AE6/r5ptTp6EPT13NzRf0G/Ou28e4KNLQnbTaqcfNEWOx2FyUukY+Nab1N3bXGt3hJOx+Wm5ASuUG8yr8ar19oJO6uYxhsqxZFOf42i0lm90fJgCt
4NP+pNr/m/2FRYLQjH8Y5cqIJtEmvYeBjKtfeWMCbYjcRWtkbkE2Id3ImEB7qTqtY8wB3vUb08xkGoCdIkSI5ovesXyUnjPxIT7A8gOTdiacLtn8Q76kK3kAF9yjJ8PM
Fawaq37EKLbP9m9woY+tXCwrqBu9pCechBqAjPC9RpEQeqfsA5KJa9abEKu+vDNH53TGWX1g24cjmT22o2vypZHDYAMPsMpX4ClOtEMmtg76tsF/7iPUDmzU1BumDRtr
wSiKNRrHB5b4MngJUMxuIMqIJtEmvYeBjKtfeWMCbYgscjoNBMu1CLtqI8qHDyz5UpEJcA+JoTc5gSn25PctGMci0tAXuZkPLOfXt1toRnj15QzDmy9CkTIbI8PjPXBA
wnhpVTvwwoJr/ftGExDiEx297J3u0rmcogtdeZMhKqGShFEPum5NWjpCgqaDqsAB07Bkgn7G+x7ZAyC5f7gbKiASRp/Sw0WzzhKwUf3xMqZHbE8R0jHvFGkRAPbPyPGB
neEVGyJd6P2vLC1LhGibNqkAGTTW78BlWWjz26dXTzeLtGD9syEqssNvAVeIZSZsHOpPxyE9MP15Hzs062pwj62WPl3UpB+JWOqJkkljU1c+jLMCkituMts2u+u0Yf9y
DaoT8A/UVctujU264+XwRZzIB04B69zUn8aMC4mxTf4eZwTMC0/rBJXC5QKs6vNwKbShjC5e+MAANF9VSB1dTcPT7bfN28N6LlEUPuqiztTr9QliMbsPyXTua37EKl8h
tc46pAiTuGC+Au0ukC44yMqIJtEmvYeBjKtfeWMCbYg5t22Fs99BiOU2t8IuD6yxlooOTciuwr1b44CPRR0qhS8o5huawvNICBwABGu4Pr5mUTvESfkktGd7xXwJGbGt
UaLwr5BdD5vS5yulP3+e0/MltpseCpJMXo1qttFjJBHjUWd8J5mQUmZonBqVVrmEq42rhFAFnzK9Np3ffOnb7nkKHMN7iXjAxbEgbUTKeHZlypYJrhwkigoHUEWeZQBK
82pQBsZ9Q/Gp0v12IrBxzeHXKSMEyZQ/3zb6MLQE1qU76/OsxPHvzgrVBUec+yTpyogm0Sa9h4GMq195YwJtiOUcDTePPiObZdx4I93XaqvygPKn2HO4TlbX/Y3GGKQA
yERaGp2S2i2zA46pdBcLQVkmSHmDGP1WUFissK36anJRovCvkF0Pm9LnK6U/f57ThUtIydkzcN1BcNquaPYIGQ2qE/AP1FXLbo1NuuPl8EU5/fov8sQ3oUbkgDvL1WmP
UpEJcA+JoTc5gSn25PctGGtfQXerXxA/M5ycVy88thC8MVflD7jjhDGQAhRgZrVmrZY+XdSkH4lY6omSSWNTVyclj4pODaFQ2o2JUvcYhwxEx7SDuyF0S5IAc1wGiFcJ
AT7aWOQwJWEU5YDL3FPAcx5nBMwLT+sElcLlAqzq83D64kLHFw1ZvG4ABYRyadsBVrwIalSidb+cns0hf2g7ACDhuFtWhU1HyXn62aH2pxbAbOZrwllk0WdgRIpS85eD
yogm0Sa9h4GMq195YwJtiNeRMuNMtb41wr5GCoDMzKAeZwTMC0/rBJXC5QKs6vNwK7gnD6h9O79dKLJ2lvRiqhHWYVJyQ0xQehxB/+UUWNStlj5d1KQfiVjqiZJJY1NX
yr15Zl+4uOKa8KmpFX7UKsqIJtEmvYeBjKtfeWMCbYioufbdq301ED3DHhUIOWpaAy0zeDNLArqeBcNr+ImJl8bInWbCFjEtlGtVsJMh2ogP8svrLyVJCsxmcUZzdvEt
rZY+XdSkH4lY6omSSWNTV/YmAn7vJ1FVU39j7VT2VRVEx7SDuyF0S5IAc1wGiFcJi/6rHTalKKm4SVIC0adoAR5nBMwLT+sElcLlAqzq83Dacw6T4dNGtZydpUJyxg30
VIOEnhIYY1XCvSD0xKNvFyDhuFtWhU1HyXn62aH2pxYU0vQ4TkQrWzwfjYVdjw6ryogm0Sa9h4GMq195YwJtiJth2LkRd34ryx6fGyZEDAMeZwTMC0/rBJXC5QKs6vNw
HTYNA9l4MxMSAyET+petKBRcSOYug7hRPJyYxKbDNMytlj5d1KQfiVjqiZJJY1NXIwh/W09XkyxUAKqg7dRBGsqIJtEmvYeBjKtfeWMCbYi3IH8hryoRzBIBYpyjs/RY
Ay0zeDNLArqeBcNr+ImJl5HYF+k2FcmdqHTmLyshxqITen0klxzc6vFece9yuGHZrZY+XdSkH4lY6omSSWNTV7Or8IYW6lT2564Eu/twojFEx7SDuyF0S5IAc1wGiFcJ
8fwpUqrCSmoSKEMo/P++vh5nBMwLT+sElcLlAqzq83AsOlixPe9HNikwkSt4xqksqIV5EW7NkRZfer1DZ/dL+CDhuFtWhU1HyXn62aH2pxa3NqyrTzzxbX1iE/uTFVSr
yogm0Sa9h4GMq195YwJtiAZSGWgYuJRv2A4lckluMP4eZwTMC0/rBJXC5QKs6vNwacbHFGpCPNmSiBMqxM8Z2Z0BjebR3oenOc9ON/hW4eutlj5d1KQfiVjqiZJJY1NX
TLN/NdrorDac13IFBmZHhcqIJtEmvYeBjKtfeWMCbYitXqmFXyHHOr9YEUwZyOznAy0zeDNLArqeBcNr+ImJl+X5E5pTPYXRNXIDVWWpWYntcz21LpD28dPqdcIfJDMu
rZY+XdSkH4lY6omSSWNTV0N5Fg3AvTHzwR8Ov82a1sJEx7SDuyF0S5IAc1wGiFcJWfOK6HSSOF972HTUlFyUBAMtM3gzSwK6ngXDa/iJiZe4UMerwfKMuKH1SmCt+BQg
v13/ZF1Giu9z/Rn+fCNRlu9QRXlbAOythLHbWs3xco0OaqneUktMxrVnWeP2ey5ERMe0g7shdEuSAHNcBohXCQhKCt8WtCk18Sq9PxvyxJ0DLTN4M0sCup4Fw2v4iYmX
+ilB02QmR5uoXMZ5qns7sXUpjPGb6kOfQWP5gxEeIdDvUEV5WwDsrYSx21rN8XKNr9z2dSfCqb75iV2JiPfavETHtIO7IXRLkgBzXAaIVwnMvwNV6ocgzOqwjgQkGTTi
Ay0zeDNLArqeBcNr+ImJl9L0CYvAe8Ve1Yiz5bhsEBCm8Ae3ovBO6QrfIH6DzMbw71BFeVsA7K2EsdtazfFyjap+YUIsB+j+f6lw1C1LbhlEx7SDuyF0S5IAc1wGiFcJ
4QHTH9DUeUYkd5MjnaEhxQMtM3gzSwK6ngXDa/iJiZdag7XTXEy/TGIg42miptM/OozK1PWhb13huL68zq4WGVGi8K+QXQ+b0ucrpT9/ntPE9ACs6igwiuG5yU37KCiL
yogm0Sa9h4GMq195YwJtiAmj5PCRmbJ/iF4fr8Tvb6MeZwTMC0/rBJXC5QKs6vNwl9nKk1f936qFiMfnDt6DSvnpTPW8kgZ2wxb2LQ/jhqVRovCvkF0Pm9LnK6U/f57T
PFWHc/jeqSkXmmgg4L3NF8qIJtEmvYeBjKtfeWMCbYh4xbzHeKAe238qAytYn/P8HmcEzAtP6wSVwuUCrOrzcBXVd9t32QsNs46pdYG7/AoEbqF7P8RO41ZVy/pCTM/N
UaLwr5BdD5vS5yulP3+e026EnViA0xwSFnm/1Tx3HxXKiCbRJr2HgYyrX3ljAm2IMeDMBb/y6+9YHriLaBBFgR5nBMwLT+sElcLlAqzq83Be382FeCz+kAQ8him2itQO
+8l6pL6YkQCiw+qwczS7HK2WPl3UpB+JWOqJkkljU1drENnos2zu/xiEq1T0ultq3tg36JZIjTN8D7VQ9R/VstViExtU/YmuwRMEvhQAPXnj2KSvYoMebAYY6iiN7r3P
7l9SXZyEhwSDyW5sMSs/Us3bNu0gJLss+nJjcYhLwlct6cOEQH9+7ZEUvNQWUJB7Bj2IVr4vzOEeL2JI8zKdW5DdT2rcUC5+gEQ/BhhH+/WHQQwKzfSgNvDjjOXRtz0D
wnhpVTvwwoJr/ftGExDiE9HHjhfC528JtN7xP8biS00+X3Kq3Txc5KDOEyQrHfihxkZFz1h9vvwLULgfSKYp2R5nBMwLT+sElcLlAqzq83Ac/rbgpwBCJAaaVMuHe/K4
n9B3BjwsE4Vb8ZmHl5vNPSpB02C2d3hVYEehXKvG/KyGYdNdBGVHlvdtWPqNImgEkyjNbvtloOMTsWlhkUC+SluIHgTS5UaP4bHyjA/4vGjmjYZGTPpx5fHkDH12aeTG
Su69n4lPbVnPBDTF6F5p2yoMCFB+ono46v6efV+6Zf3nQEE6sS8QwG1/bethI6hcqyks6Uws+wRR+WVIcJ+QKCkV3+NFkZrlvNYQ43QWj5mq6sL5TWabc1JCcYR6AYY5
uY5z/UiHUqwsHvmOrlepRKHW93jL5+Orc7mKfNhHQNYnPUyPFVX8cKpO+ySb+a3ILA5E86rW/lPsHTKaF5kcfOPYpK9igx5sBhjqKI3uvc99YBk6vVwhClgf3ogYtSLr
zds27SAkuyz6cmNxiEvCVysCOMbyfGbwV6JN4CcNUdLenDyZZ1OcbTkmDvvGHtMpzRqFSenvVk0sY5jJJpVNhMzqLsTLB5OCqxGlycKVmVfCeGlVO/DCgmv9+0YTEOIT
c3pYleE37TbzRaUQ7BAT5swH71xp2I6eRNDSVOhy8XpbbhswebkcwWiDxtf6TUsMHmcEzAtP6wSVwuUCrOrzcAsUMTkbsIYDanN+xIxV2RxKP9upODCmAvFJm/5wCD3m
KkHTYLZ3eFVgR6Fcq8b8rOIdAoskcL9Aket27w+PJVtHbE8R0jHvFGkRAPbPyPGB6UMk4u/NX8a8cxiUvzV7C8qIJtEmvYeBjKtfeWMCbYiUMg+ZBGvdlKsEM0bso0rt
koRRD7puTVo6QoKmg6rAAQKoIJ4M3RBhnCktY+NkdUSt4gDPKy0gXN2S2jIKm89GMJCd8nLEhVrX+ujqZJgSi5Ab1eIMCc8ewPhoWmfm15Stlj5d1KQfiVjqiZJJY1NX
KyBByjOI0oo89PEgUWmkVd7YN+iWSI0zfA+1UPUf1bKXE9yviwrWoVdhr/ygGb3049ikr2KDHmwGGOooje69z5rzf9M53N9OH+85wAJlMxvN2zbtICS7LPpyY3GIS8JX
9xTRFj/rLJFGuPU+aoV4bFx8q/OXOJSIDv1m/TN3RmCQ3U9q3FAufoBEPwYYR/v1gwgDEPRTe5dUF4LOFK9UEcJ4aVU78MKCa/37RhMQ4hMnOL7MbVrVpWAOJyYoOE08
zAfvXGnYjp5E0NJU6HLxelXqLLCzLcEXOj62poMz5IseZwTMC0/rBJXC5QKs6vNwrECYEr7640IQzqP7L+HqaSP1BoreRx5yIXL3HnVZookqQdNgtnd4VWBHoVyrxvys
l/XfaBWQD13mhqc38L3ZAUdsTxHSMe8UaREA9s/I8YGJnYdOagOGg+b/DNtpc0kPyogm0Sa9h4GMq195YwJtiL2hpV45dO7oGu7HRUfXl7qShFEPum5NWjpCgqaDqsAB
JnfEUOQSuy0fI7Y1zf21eYcySvn0XPAFGsul0kHzdfUdSOA8Waq8SxDnzh76k8/MvS2D+u6R2on3AuTwm67oaa2WPl3UpB+JWOqJkkljU1fCJJTIZ11B45U+vKUG4Cb2
3tg36JZIjTN8D7VQ9R/VsjAVMz3t0nPw0dPGbbjdFG7j2KSvYoMebAYY6iiN7r3Pozx+5P3/9WZu623gLIG4Dc3bNu0gJLss+nJjcYhLwlcDTpGWC82kLioWCza3ZCXT
JzXnT741Lb5k3Hv1+7oSh5DdT2rcUC5+gEQ/BhhH+/W+OGhCvsUY/9Ve6RRWqZxawnhpVTvwwoJr/ftGExDiE6/2avET8Xv1fZJRrL8GCh3MB+9cadiOnkTQ0lTocvF6
0YLDvHheidgbjdlJiMAqYB5nBMwLT+sElcLlAqzq83AZgouTQc9URVrQUxhP+nR2cUllVJiGY7wHb9XSCzk5yjFiZ/1N++J5mriLX7iVoF7CZZ9SGx9sFNCI7prtT0gT
DT2KOrsT9gjx9wo9umnRP2T1uvRQ5rM/3NkM2HEjWi+Lkil0UJwP4VVNvOw1v37ZXem1mAkh2wYo1dPVVDH/wSoMCFB+ono46v6efV+6Zf3Uzk2FwTXylOufQbohAsM9
tJr3e48VlD+CLYF7F/GNE6FE4X4q9l4Xutb/foq2wDhoBGKix2CZ9qLg2tWmCVO4uY5z/UiHUqwsHvmOrlepRBtw0hvjo8e29tj1Otbx1lvSTGeObs7fK9H/zE6InBQ5
/8K9jOmdsh958y0WCZ0FSAjNjxZSbDLkWIYr2E/C8jgjG/MpOC5Ocl8LY5rTpJqpgYEsXK3n47fHF/xXpmDOs16il+3z8jc1VyMaIWpDL5nQ52nJaoJDWd6Mr/T+Lnen
knVfFikngIHMkgsguEwexyFqK7p7IRdTDXNlfQprozBPij7JwWM0tqL57l8VlYPPYhVMvsNNK4PZY7FBrYoUlMqIJtEmvYeBjKtfeWMCbYgmj2IFBQi0L2hjqjEYsUAe
ylDCQKCml7o7S7hDp0qAIK2WPl3UpB+JWOqJkkljU1dcw4SQl4zT/JeGgsyPzzsuJqb+RVARH5TYV84Dt01m8B90bT7nAzDZAZdiyeeDUaQZNqmrhr6BvfmBg0OjA6V6
Si1RC8IM23su3CdYkV6fBvyywkYVd8nfbEq+AjBGRbH3y1kNltoKNxBZqT/K8DCU9BIBnjz+ivfNfGBxGhHcyOH/YZ37gRlU1xjT0kRK2jQa8lI+zLPzyF2wLE7YZVbl
L3Yi4mezW3hmn2I1iLEkSXG6Ez2CnIRNHah2w7We/hDEZaKtK87dtq3QuZ/fySmfc75K9hEEpxZ9vv8oVCUpahudnWZpo9leaNOjc8l/HsdfCkARKMFQ7ZfmzOgyrVHn
M45f9yjY3jTBMWvo6TdXvTGWl2qVXUaqe3X+h3ll45Y1XsJa63rNjsoWIXyOjZ+mj1Q8h+53WwsxPhI7McAhNyL+WGcI4lxDo2hbK8G7IJtHhFHI63rZUmqif0+Pyh2V
GMaeRSyAzo2AEa73z25Nrou4w+YVF7RY4CjIE0+WvzMcTgF3N6yOuiVrUrYgVHrScps4xFwK84996QooV3yQrcfeplROp5QhwSa9stUG9QblSA1zKzNZXa+bey389pNd
5NsgWxSpbWHTB55I949rgmw4YIZ9fuybmueYIRikK15iXwSqpNOfH4lj8DuGxmQQk4O9sq9hu3LMciKcudDkVCMxlr3fI7eTX3H2wbR3fLVOn55EZlmnRR+6WV3z3iwk
tqBgj+1AyQvqv7HExQUlYQ9WR4RV2/X1sw0p7N+HaWzwSSM9Ox6k4qEA9cu4xf3xDW3iry758mTmz8eX70BaiEq94N7QY6UEFeEuGm85xxprIKydQN0/m+Yqq/YKy+ul
fiaj/1OM91k8R84eCwE1OMMjJb5EJpdo3xVAR7F3mlL9w5Gwv76d82EwCnKeOwrjXDIhnBy5TEwh8TtfDv4ZpnnIuZ/WFMqPYfIGSIbbO14H4kxgaklpAo734b4yeNwj
jRxuJB+8fmyLTzcR8ONlQ7ac7MX0YFQB9C70AlP0sddYzxgEZYD4P9/4yXFVBBtO70TCfwzyXSFw4BkAoVB1Wr8w/L/TyAHl6ya5avHDve4zTHwCfWRG408mCWP0CV5T
hlbAETp19o2p+16W3+IUNhku9JBx95CzeGbnL0MZ628bFt9dq8c6ReF+d+oc7ZMqTe8OGoy1kqP5CD9DquzESFxYlkG+Ok4lnjsW6R31SS4iLmTRLzhXplLyo4Bcw3lV
uhBqKBnIs1+C+yMRYJSmVPMskxaJufkU2PtMup8JrNfLpK3sKcSvezoVff5r3+M1gAzVMq6U0ohMe+3O6QYJJlFA7VdhtWq5pARfkaMssoKOEfMyYXt5HPmQF3upyAS2
1kSHWwp7wbu/6JsZXxGqb0Xsgo50/S7EZNb74JzJYyEz/DLipR/okN4KGMbBtR7tjACU/N9e3ZgH7KoS65+hbb+VCzpbfEAaFX7dYj9tmGZZja+AwrlxGlHPV8APaQnZ
U6bgO2hzpVM70iDAxRsbW8UpV4/EkMTFdHjLeZsJFAjLpK3sKcSvezoVff5r3+M1gAzVMq6U0ohMe+3O6QYJJg4YV/NOG5nFs13Sb61xWztTBmoWuZy0yJa+iGXEQZ9F
DiZSJpmOWZyUxjLzB4HqzESuqtFaC4ssy+ITOZpmGMe/l7nlr/mlcamM+8eW2AUe70TCfwzyXSFw4BkAoVB1Wo+CNshuZ4cQm92PSFNkI4DstaQH54KvV5wS0KRjA3vz
loPWl4j8R4R4mB6bqLENPNchdOHU/fp+Zqxg54D48QQrZfFcd6iJtel2KERb6d8IZJq5m5zK0lss1cSNcw/wyI0MXsywLPH1jMspHK0EgHcoPr61vcRYZq7x3rRhVWSO
7C3KpEcCZ/A/f1Sil67zQ1cy/Z6R2FK0dLPAmhvqUmkLflRzsV/BzXEFNb6L1XDihHK9dr4rOrY8ORTHfJjVtO0Bva8ZomWPX8rQjF/WqTA2JBYM7kHKWfibfkO5nmuZ
gzCV7Pu5vCEaXc31VByhXQtV0miOmsB9Q4+4f7jA3Ri9gOjOueFcFyN6nT25c/LsmjLgQBgRAdsXjhpzErIo81A7o/QV+LluECImEpMvD74+mIQSFz1raxKu0b9je8vH
4G5Bgeua26Cp2323v+AlJrRlqvnOhCW42G3yfmkP4MwOQSonnyZJLWKpUupgzNe63BQ87h5Bit0iFYpo+xeEYOdWdp1AzV1rdoSslZ88oGF4GbOK5ik2bQJ7mDlBgyxB
5yIM9OdllrMKvacu7WJvC+NLcGJ/LNlxGntA4oHaRzF4HKjMN9dxHnUhiQgNBIIk2nYSqR0fMxsYG/Hgu38zaYo68NSyMRMXatl7LfdP3K3uG6Q/OWypj4r2wyyXyJCM
0DsOKfO/hSTCcRQ6HkLvOoNGeVNUKb+VKlqDGNZNG7rvRMJ/DPJdIXDgGQChUHVa/oUzK7Zwww/1yjffScUD/CK8S9DJhrnHLVXqSpEGkOauWktFFNsQhmwL2Cb6N+Dx
bF82JbVLSZYq0fcHKVOiSlW1RSytyEkPvyW9FRZctC6STKcYjofvHyr6qf2GdtEnObVLPW2ylQETyXZCmphdNno+0oEeZ94n1Xu6/+00jR+TvpQgS+8MME0frzLXZ4LZ
C1XSaI6awH1Dj7h/uMDdGOdup7wlB1Q5HAYczYIkFTaZzGUXApFtsSsfWEbgr6oUWER39YYBlgL19HkXxBkNPvSg3bEQVKZQRynAAyGZi1Gg2ZK52vF6uhejEnT/XXcp
JGT4Byu8gAAEHU9ABcUOhRIXHJcOZtRWAFoRsUHJAcirsx2gD5hxoJyty0eoPKRGKA7x+SaMKUbwmHPdx2zd8rFtjzck7+TxES1IMamTb/DeNgbyazXVi61v6qLFuiik
ZtMkRI4iXSQf3xR/WsAdw/IyngSoc3LXW9fb+fijEQSaHgPfNnScwJ+yb3vp8eFfdZS8FfD+3GvAhl4yggUrCz4pwIIj0NC5exRonTpd5Ifb34VnHE7vFMukW0S2HoW4
XuliOb4u6YIDMKyJJjwh4+MozG8Ghdz+vATtTWUYErRlWcUUM/dyV0+rGiAJG3PZKhLpWKyCnFm3HUvQljioJCv6wxOyLoohfu7gxOhas2+cG9c+NP0Z6To57WrqCIh7
eHb+04VcZyvvPAB1WxhB9+a4p4HlnMmFRM5jWRcGiSK/v5aQ19LdEHYhHVKTTNzWl8PTD59PGw3bYez+FBSCUPPYtOyH3DtF4l9lY/9ZiWgmQzHiyeSHOHxaOsZQf/5A
SwOofqZG8UkhGwNh2rTmvOsUGkTI8mSSdcFAq4MATLab48h1T9+6cAuTtt+pcD6bhSe2ZfPgRTddKsnkPP7IgGXukBiuh+3Mtss7hLjaziT6jwntKAW5KiZgF6r1fDcT
t2kAuA85O+gpDP8RVfHFyZbptWjmTQFlpMrjJMcaA6X31wb4uNO4WMfvO3wJZKQKGKvQ36ed/njFyl1ZVYesR9vfhWccTu8Uy6RbRLYehbiGnuABIDTzzQzpK14XFqhX
rfkrh+KprEQsNP1uS8QMjuLdET0teE5ZuKn53e6mnl2gkbv1C3vmctIlMTWiMRsu92TvwYkIX7UC/NT81WJP6Cv0j2on4X8yDfQEGfZpcP1Ah1P2iA6XBkTDhnca4F5r
C1JePAw3HHZjoxtd7+9GC1d/nUQVTj1PQfXmrM6cPmsj5k1RThuDQsNbndID4MM2lxL26b911tryMnrWPXpBWcOYOdb5Qw1sGoSu2Vn+jEEXW5tgBD9op3MqbgF0up4t
3zN27xT9AGNUNc0RM9L+cJUe0InaU0cZDx424g50I3kknaehv1pULqonS+ZGKOC2VVV0YJ5crQnjgGDzQsLyF714ji/Q3WFaGIkwxwyLEyG4BVn6Eb/FrCrZGp5fZmKh
Ij6EcV0AEM18TzI5qwyhw+TYprblJBWlgl7IPmmhnq1Xf51EFU49T0H15qzOnD5r4SlJQTDy5MeIgqw/alDaNZcS9um/ddba8jJ61j16QVnV2PmYkbvUMKP79CBMpMtR
gfvBwCQvrBbAYt9N+FUbC7EIJwZSeoHfUAHLI4y2Fhsze2OTxf3j7aI38C9UNHvqEhTVRaUCF3er0KOVSMIpGUE3i3z03CxGWHxjOW4HM54gE1Slu5rQDGHN8s49p5D4
LnBPLbCjOLf5W48WzrdlR56NVD9nV5pW1qbVr6SyGLc9gfzwQk51BOLTcq0FGqfWZk++MkJ5mSpLNq5rudSuou1uJE+z1tOsSfXuN5xiemaLEZOUQ1wLWn/aoy2oCdFP
KS53Gvrvg0nqUuimtVdC7KPJzQDWJKzSmegg9bYI2YU2ItMGMHVL7EKzqZZz8K7pjYX4XLjun2wh3SsX57xk84wh9s1ez1whMgjCok7SqIqQvChoybHUYICKt0hkdgnl
e8aglDVaJR29WmNJv6ePi6C7kO6xwwG12bO56Z5eL15mT74yQnmZKks2rmu51K6ikKxQe0HXsEtTdPWRyOcmcIsRk5RDXAtaf9qjLagJ0U8pLnca+u+DSepS6Ka1V0Ls
UdxDHm4RSWIWVrb1UIWn4TYi0wYwdUvsQrOplnPwrumNhfhcuO6fbCHdKxfnvGTzaG4QNtM+uYpaOIITUTpY+ZC8KGjJsdRggIq3SGR2CeV7xqCUNVolHb1aY0m/p4+L
NvUZ8UZBy5sbqK4GHIwjEmZPvjJCeZkqSzaua7nUrqKvnXZbsO/WQ5erieUffUTeYhbslfK12de8qZ7ws3Y9W/gCIhcnluy92at3eH0oox4ucE8tsKM4t/lbjxbOt2VH
mtAvo2TtQf6v79K0bGY1VRRQl62+9cr36jtaVM41fVcpLnca+u+DSepS6Ka1V0LsVE0nD/sV/GS+OXVg3yYK/fFW3GQQPsIZMahHCH1ZfwdntSGW27Gz/mRkarbIB3BH
CeCFZQaFBsAVc7nn5ATq5aD7iN1Dox7z56JbGvuQCFo4s1wFkJ5VPIZOm7N13Qzz76OJPV6T66eL8YT448mD2zvtDHXdZZPhr/y9MewweBisapPODQ3Mq2OTIWlrX36z
GlH309IX7eqMTCJXF1ZxY/ua2mrnQg8wwr5snmLrwpg83ja9mTJudWCmlMLGQGruSUfDtNGWy7noAQpT0MVRLza+AmcSjCjH6Mk2L83HbScpLnca+u+DSepS6Ka1V0Ls
Ky2/YTtV0Nj6S6zoSOBhPwSv5eRdVmPY8dPgzIxjdyX7mtpq50IPMMK+bJ5i68KY2b0DW70l9DpNHe9usBu1jtebV3Db63+n8Yy4CUnBy58J4IVlBoUGwBVzuefkBOrl
F/nzpHBZLZxa+GHvktK/qREWsJ6lee7o8V88xF5RGWvtnWdliBzyQNEDHQhf14L87XSTFInTTmAK4IlOx3M5/tcclNgaevUsdm7dIZQaRdyNhfhcuO6fbCHdKxfnvGTz
tyGZHAlrcTagBOpOT5Xr4fn1XbxOGQ7hTjMgOs5xF/+FziNLDMOyrZbx++vwUaAq9saXafw+LhZEr8SPz4yb7z2Hrx9Q4Co0q6/2U8FGzeUc+6HMlmOsQQUNo1FrCj+0
n9nnyQY1z6WVccJHKrBVtpUHrCQ+kDUcSWo9qgrOKisucE8tsKM4t/lbjxbOt2VHxBJ1zNy71unevzWuvXWxCtxO1f+DJ1ugNVGT8HM3KHF7xqCUNVolHb1aY0m/p4+L
c2KBfHqLC7U81a0bgI85Di0pP8K60AWgvOM4TqIUuVwpLnca+u+DSepS6Ka1V0Ls8Tt9AqPYs4Jxa/KTPtc3s8vQUZdLELwQGB76c30AzTWSNKX/0s9NEKY4KNhQHnlo
jvfNrUD13fj5IvTImmUKV6wWVpYgxIUhEJZ3l/6hE+hHeN0Z9fFVfh1iu8WBxXEmyogm0Sa9h4GMq195YwJtiDdv66OnVRJAau0dxUGai1vKiCbRJr2HgYyrX3ljAm2I
KbAWmvuvd8ilV1icDV9dy6Si6wmrysR4iCuu2qvqEoTKiCbRJr2HgYyrX3ljAm2I45UR6ZE1bSDQ1wubuNrH28qIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFG
0D8ArNmKT5z6JR/X5ZWW7MqIJtEmvYeBjKtfeWMCbYiCX712GIgul2ek6aITwKPIgcrPEumJRM3yGBMVWpjK2XIHLql8/FShcQ41SVHzY3bjuS03TTiHdwe0LOIJRTaz
yogm0Sa9h4GMq195YwJtiCjMrfZC18kZgmyexZprnpDMEOrDFGST6DOvm+tIGKSJ3gRHoQ0bubQUMPVuAEVMOlZDNNcbEKu2GTB2kCKnikUkx3bMZuA5jd0dNaF4flX9
UNp1bqmHVvy30bZRA1z2/25ePDzMcisObgzj5ZFSfd/IhhD76vmdN72p1ECVhN29g5EujPTMy563mg9xoD0cXcy++cnVCkCopZ9VlzBXBglJld1HA3ixoQP+zzXD+t1M
BL+P3z60IV38x1jPgNNd+jTER5laSx7c5M9idLzk32T2uzAflGXdSR4nP5/retPvjkJ+lfbPp/2c+EO3keUV6MqIJtEmvYeBjKtfeWMCbYi9Ovw+7QQGVJKO8dvFnQoo
yDIGwD6ItGTZtJu2QbM0YenHVftzjYQ56eym/QM73ELP8hujN87nCKzCfCSbGQkYymm/k7uRFFpLpKX9AwZ0CGsikNY0oYBf0zpBRx2Hwp844Emp1nvdKOlkxC+0i3BD
SYzVIdJIh+US8B5kR7PJB8Ya7J+CiiRRsYsnvbOEJyfRWKSqc5EX+h0bd7wNrMhnvKcbwrKV4pP1PTyOXXOUtRGXK+pTALQuvKskpm39surLpRlnVr7k6QshsnsuR6lA
wBqJVfqn/L4hfdyIqDTh15dJo1EWvLurCBlGuyDlBw2uyJU+BiEPWy05AZ+Wr7d4OOPxh4OVLHo6tCilgvacitN4D+wHk19YOJEoBAac+tU9jZwXBfvMF8OadfGHNkcW
X0l1T2q8lxvuQs3gQl1nD8kKh+D3K3YJSN8zpkS7pT6LMtawqsVo5gs3KrDV0oapDGn/Ut81LfZoWSUG+m6lTtL2fwuQ+LsVfIRkdOsgMXPyspLUWNhXIn5bdmxIBgdt
yogm0Sa9h4GMq195YwJtiKvhyO7aWZXkK94E9Qlai+yodW+LnoxK82EvIPpOAfXhVojj5TLzk0D/SFDJrfxWCZadnmUUF9tCzXGoZ+EtNU/KiCbRJr2HgYyrX3ljAm2I
XBYojzkHB78N/tNAlJgvWsqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iq4QROTE8Ou5/BD682au49m78WJ7owZFWNE9tsFuB5ZbmXpFp3HejhipdKDgxGKw1C
FXlkhpt3pfqPbksifPqRHTRYlTE78nku/iN2dKkUNF+0VwsCiyKmkiqkVEPh3bRLagCn9gkK7gpLgbxgv7tce6gcPGV4pFAmbi2MlKQ4r5+8PfWzYMep7b2QLXWXV6xy
yogm0Sa9h4GMq195YwJtiIaalFuVVmXMEPxu9ZqMuUpBCaBDS5gzAmNw11HlqrYbgRrInBgZD19HN9j5BZzno/VGIlHRJYcLy0uwOS+262KxUpBEHIYNAgisGtBZb5zq
NzbBk5wDw6YZhjQ+XAyYnG6b6XIrcUR5Dk4VMf5tb6101vl16HpxIuZMEoNeozDPHzMgG/AjQ2U9LqcwqzUbbSG8E+/izOgDZtCcT6SY28S8pxvCspXik/U9PI5dc5S1
a4lMOuQbvCfDrDUj+m35aktFicG7TD+R/KGPyE32lKJWQzTXGxCrthkwdpAip4pF9SWHxLlJdJ2AVUfW6nvva1DadW6ph1b8t9G2UQNc9v9uXjw8zHIrDm4M4+WRUn3f
vlm1ZWEZYM0ySa19UwrZYffCP/TXf2t2gojDevOlUhNJU+A8/2h02YhPD1qTo7H1yogm0Sa9h4GMq195YwJtiIaalFuVVmXMEPxu9ZqMuUrxw5NVMe8YCiXOiyFM5vQZ
fUgoSjZJ0mfLOvTfraoVzlffkEP7Y9sZtTpdtZ1RijOxUpBEHIYNAgisGtBZb5zqNzbBk5wDw6YZhjQ+XAyYnCayXQosBNtXJl2WW77ohEB01vl16HpxIuZMEoNeozDP
hNfsImzUUfGrOJHCGDefGYanyWygkFx8mtgge9EO3CO8pxvCspXik/U9PI5dc5S1EZcr6lMAtC68qySmbf2y6kh7E8ibURM9QIkmd+eOIRDiSUf02i//vvXpnXzJnRhp
xEFWkkRPRnFv/j0lZ6r/nVDadW6ph1b8t9G2UQNc9v9uXjw8zHIrDm4M4+WRUn3f2pgRUJvbeeSYtIpd3p3A3KmqpWVKVlD55lizL+l5rJBszLK40/MhgE/ai76XOxxk
yogm0Sa9h4GMq195YwJtiIQBQ3d4Eg+do7dTRpvk0D7OgNn+h0jGzwupwl3UCMEpfUgoSjZJ0mfLOvTfraoVzjGzhEPTiwRKqgoj1bJ3VHfKiCbRJr2HgYyrX3ljAm2I
FOkkgAvTE+UMiwy3mhb1lwCkaqtri+07+j4KEdNZHBN01vl16HpxIuZMEoNeozDPXOeR5zTyZnOOQfinxhoykf2WBQ6Ad8OImCJ/aGgwP528pxvCspXik/U9PI5dc5S1
EwHQn/r7znhvgyNwTVDexgyDVHNcft/H/V8j6QDvPenMLUdzy1MBeF977l1E8SkspRnVJPGydfTNfOffJx75plDadW6ph1b8t9G2UQNc9v8eA+DWbCA8EOqFHBG5AnJx
X88wVpug7x6aqRbU7fsCL6mqpWVKVlD55lizL+l5rJBGgJovLVwVoD+4/Reh5e2Gyogm0Sa9h4GMq195YwJtiIQBQ3d4Eg+do7dTRpvk0D4AcKb/Di1FW2zkdyWXfGHz
fUgoSjZJ0mfLOvTfraoVzslE0iOX/2AljmklfmnssHfKiCbRJr2HgYyrX3ljAm2INzbBk5wDw6YZhjQ+XAyYnFzGdVjkvlMGAdkQI4OW+/+N3JATQDmfYCyLC0DOLr5N
9GQgm3xOhDMrU9WYsdJKeItga29j9WzWHanK0tEH3sRqb5eRcMom5Z+FQBdfyjYnyogm0Sa9h4GMq195YwJtiN4ER6ENG7m0FDD1bgBFTDqxuQf9ZvwJc/2CSs8YMsdP
2MZjK+n+YhsmZ81VFDwNMKwjK3BzueTz55ezm5Vm7pOC4CrsfS0J3Ue8tl2Wmivm2pgRUJvbeeSYtIpd3p3A3CPyA0o2okRxHprUNUy1db+9rENtjWJHQ229BSfCYqYs
yogm0Sa9h4GMq195YwJtiP4/4w42v55BjTY1Lh2obofKiCbRJr2HgYyrX3ljAm2IgRrInBgZD19HN9j5BZzno6nDPBcOr/9Bnx4cY/pv35hugE88QuHUpugyFK4YQzL2
NLTk8fihr5NpSyt35tv0ty+VdF67+03VgYK29kzvLJB+yGZrmBneblZRmw9FMfTX71KPw0RIXgLV6qRy+WoELTa98/mrWNaN0UqTe9AiClVRcmr3O2O1bg5FOB5w8dq+
k1vLDD1jj6Q+n+aRuddo2I7iQ7nBaKh+iDx0aaXgHgAxsUfkMkvKO8mmX6YN8HXiBobYEQ+Nh06EWNOfSwHiY5bAFkRIlETukh5yM2ca77tU6co60/5xo+OxKJHfFKod
Qt740ybFOyn1xxQWFfZN1fDuFpFTYUg8RVN19ERnN4vSBoqsTXZBfKS4CqWNm/178xXIL3kuNLnW4kvgxoGJ+2Ig0J81fTpbl1WUQyKhaRQV0mRPfb2LsI6eEzUpjEqh
X5jNwbBY5EShrOd8GEjjtSqPZvSsJfn1fRBz/Evb+4rkitwaGdT73c2EeXEwimmyCzA1giAT9fiKUkIvtLOxqq6HwZ8L58XqpY/cUSRxconS9n8LkPi7FXyEZHTrIDFz
mbKUgndlvXpXTBnaqNhCwUmV3UcDeLGhA/7PNcP63Ux0AWMhoy32ZacoiagmR7C1yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
5o4oKz3coinVeeRBFcqO/nHppJYjgpGkgXvbawejv+///XTWyDbRbI+4bxUuBetlyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
RDnjCNXP+UwP9nlgWpEM3aJ3SiBZNStaEB5FbOxR1/RJtbgU+uAcoZXR8mGuIlTVbTGiGNLNGzy2EsRf7D6gf/jsIM+o2hQ63BcPX8EFrISBGsicGBkPX0c32PkFnOej
GzN7WCWm5VIt0YqQlAuoZvf0FAP1fkXsAdvbODmjCdCVZj0X4L+EhLl/yPPVTYjiNLE8UnNxW/iUDAHQJ46PyWonQ744EuFTVFTZQS9NLrwHiB/b6e0wYMey9h6BR8i9
0WlqFqBWBr1LOBmWT3ZE2UbDBD2Gaydm7eCJf6FJCx8+M1n80g30OL9EabcxTpXvyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFG
HaDv9Fo2BT80j14LCBWwtaV+Hqna1ikhIA50dr+P6wZ8mIsN0PqNPviVNLV6PE+8yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iq
h2uBK7gC6QIBLDLw6LWsc6378hrM6nGISQO8of0zsurL4o8/2IkGAXivjsMiLlEGHtJLa4LCBk/QpJrL5CdRIVloL0SszRVtItgg/Jpeay8dVA2dwaDGqbqPPttUrcNb
hs+HEGL3fZ2Wy7qYGGC0R2C6bZyR82qXuoz/t8+TMR/dOAUDVRhPk78VWoxKDOx5Ms6Yp83sbEijSPVFltsRMMqIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N2
RPSVlqBUKpiz/b3JoD4gIK4m5bsKIEjVOIq8zWedUnGEyFsz2zRis/dociCaomz9AuocZcRiEJ9sgcbvLV3atlg0UampgNzi+7SMYVfw6lMaUlSVVJOGciBZGBR8XQfQ
80s1u2OqHYTm0Fd/2Mp/6H8A/j75oRxgM/gBLozR09rbEpVtaCVW+z9C6bkCWoC2OkVpX1mPJbS8oIVeXeAfbx/1IF9go+/3/s9uyYOry45aDDdoNf2EBmp0ULiveLwK
eZeLRwEE3MinVTuLvmGoIAyf5XeP2YbbLk8URqdXMJFA24bVgXQMxBqg+LqBsqdysNzzuRNBnsXJuVOgboO8mpcKBHhjfFtwMzdJuGYXGe9qrV99K6Buhhy2PC9BzyTT
3A/HQUAYHGYwc9euKnMf/GfLqyCudIuraj9d/gNQA0VtmhmbSQFu/4QZ3IQgMYQ4tpzsxfRgVAH0LvQCU/Sx10DHmBvdcBNWM4eF2aCsD0oy4cZoWKoLRVrjQc52GLJL
bhPCaJgHQmhd4PWX/OFIGW1ZeX7aRwMqzlB+HxP1ozTkInEXnwPC4/4rNc3ldMDDyHfX90Etu+C/RxWSmaPQ8vnmzcXYi9xLwvLlzYY8oE0Xg17f+0FJ2HrRy08/29s1
bcx9A3euJafUPZh7l1vZhbUr4xUHcTLKX/ySCND/gs6O4kO5wWiofog8dGml4B4AMbFH5DJLyjvJpl+mDfB14sCd3b84K5sCXKusIxcsYqquseeuN8/IQ5kfT4T6q8t6
VOnKOtP+caPjsSiR3xSqHTlpv/7rMHRZWxzH2xuiX3nw7haRU2FIPEVTdfREZzeLnV+Vuyc4u1odPJAoAM2c6llY5rgea9KyOtkQSzEckV7XJ4ps8BDtBhJsiekfumSS
dEMpVk0/iVLB/Xc8gKO+A6qo8kgK0QTqrGTuile8vfIqj2b0rCX59X0Qc/xL2/uKPTCOW0L6tA0RU/Uqf982LqkQQwyrnNy3L9/n1qdgrTrafCmsSMQn8ESST2WieBIp
ql1NB7U/njFU5faCQY2X1+1BFIfeKwXapivPnCzKL9hJld1HA3ixoQP+zzXD+t1MComuWhI0/TMUIsz3abcxAIfPnUocYhLdJQeboMcSy2lI9QtcGHwySfxMBlCost0s
9rswH5Rl3UkeJz+f63rT75H9wEzooq+fUsQw3xpXFpgc+TaNxDDi/A0Bd7t7rbQAUMgCsOdd3THJRr23GJArZwmqoggm2wf1OP9KsYqEGRskhQiuwNeOpuEhYZfmjh30
OK8p0jZCjvddAT9CCzxkB5dP5V0IOVKk5YHDlijqBa3Qx2hjW1mZaISm6tkpPeuGgnVXWJdrlpoWPt54kYLtFg5pQuUrhjkblzQeOns6JP5c2yG6y5Jg/Bf9y0dtvLiG
biNtkv8ZosD41nbzsqiysJXenIloMZ0l4vYwk52Rbmz7rICpy6vrQuFpgCGDT3b1siM8eP7C5UP+R8TDmT/lHf9aPE9sH7MI42fPI4d1a3kjrI9FM7ztkukC08rcnFH0
6cdV+3ONhDnp7Kb9AzvcQrxetCRT4idQs8jA3m0o/pqxUpBEHIYNAgisGtBZb5zqooQOPG3OcfrPF0EFXlE0dgi9JRYLPs8uhpFWo8kbyAITl5tNIG3ChFhbIblUPuCo
nkPELMSQBI3KYVRngPExRvKcasydWBehMi8ua/FMhg6UVNyq2AQPD9kvJB4JjOspPdhOEv+mhNckXSoYAbFWIv3DkbC/vp3zYTAKcp47CuPQAi8Ea3IOEWjfZ83zpPvb
qEG1siCVfekN2bm/gFcJo9oeFZ3iSZleDixYvPEhwK77rICpy6vrQuFpgCGDT3b1dtP9lUIO57/l3EXRUcfl/GdyQjWL9s7MOjuGNxYddafXsGtl5FAi8AC3hMHSk0WL
g3EXTn58wwiGNPL7MS7te3wuCEegFy4Sxost61XiCXSsQSJa89BJLYvt2w0TUcnM0iOvNx8yGsuBUNl6SE4EbH1FKE5fikB3n8aah826wa/tWnbFSWDv4m4c8pyWb2SA
HBBXVMwMHzBKhdVnmXJsX6GNuihNM98latsGeoB2Zkwzpu9l3dXPx7c1mv75CSFshMhbM9s0YrP3aHIgmqJs/TRi6/Q7+mjbCiqWtUGmNqzhHQtrLd+Z7cnIH7JxEP51
0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNXkfl5KZF9gbEQ+eHxe+OkP2xKVbWglVvs/Qum5AlqAttZA3k0EnrdhFInzGNbJ/NwdiIojrXJTEu1goQstByaY
eMBIGBQfEV9VfZZ9LJbCaDwTKEgPkf+G3npp/y9Z6oW8ZjnbuM8AclaTwktFLzKdyy+FSkzFtYWI4MKvBJonFr88DDxyqIVgSatcicbH4t7KiCbRJr2HgYyrX3ljAm2I
3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/xu9gdMyW7TUvynp3RrYWBsbZoZm0kBbv+EGdyEIDGEOLac7MX0YFQB9C70AlP0sdd/v3C27lE7FU9m66iSzh0/
UQtKb+fYpkoggaoOn6jJ024TwmiYB0JoXeD1l/zhSBmxe+QLHCjD0Wl9TQm9f/zd5CJxF58DwuP+KzXN5XTAw5GlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKU
Gzhu9RV6EOIFkZcp3lZ92BJGqJWn1t/qGroimMFAGFbaypk9uT+rpzUCFSvQRVvIjuJDucFoqH6IPHRppeAeAP+q5nY7WBv2SyrLHBK7AUhI1mh1FNCh8htDhUnJ/pgZ
Lk97UQfGbIo8n8GY6PBTrh58cROfMe6s7K9t/3ng+cqE6xh8ZNIfXeTZ+y7XGjHk8O4WkVNhSDxFU3X0RGc3i9IGiqxNdkF8pLgKpY2b/XsGhtgRD42HToRY059LAeJj
TgT4QtMKn2r4tAPdeNFPfhXSZE99vYuwjp4TNSmMSqFrur8f9WycP8dnCGuTwUrIKo9m9Kwl+fV9EHP8S9v7ij0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4
0vjyatqlCOINRHPb7mRDpapdTQe1P54xVOX2gkGNl9fgvkp/LWqiEUPmitZhbXdfAm5HG//yPBtVhcrExLB3xKulj06rOtMbdVH1RwKTctiet466qApO6GbyADyw6Fgh
V7Sl9CKggcEMfd4nV/rtLEDJqrCQCDOrgCkmTBNGpAzOecbImhxA+FREVvp4fFk+iJPNp4FDN3PZsXyl3lw0MlDIArDnXd0xyUa9txiQK2d6XljQW/w7Z13IrwbcKGln
+QwmLyladjDGuSkGW1o9P4mvX5jRYBoyP+S0/fQvdRpjdN96IAe3AQYsi6NBFtCwxa/t7LgFOQcrkCTfih8TiYJ1V1iXa5aaFj7eeJGC7RYOaULlK4Y5G5c0Hjp7OiT+
Qk+mmEFVn2Nnda4Pf/QeQn1IKEo2SdJnyzr0362qFc5BW3ek7V/7haABuNAj3PSYz6upr3QdzVPH7b22FnMTY7IjPHj+wuVD/kfEw5k/5R3/WjxPbB+zCONnzyOHdWt5
jffVHdp/fBzRoDR4IDLJaunHVftzjYQ56eym/QM73EKiLtgP+Sx0MbomDLBjh0VF9GcaUZSFfEuJIMsRb/IZ/xNu2VDnAmvEYyiV35vU50Z1wLoUYjnAAEjwaCBgCZ6K
F91wrmGxhwihTd1JtFg7Uo9G8sc9Ts8IJ8v5APiTv42bcZupIkDSwOCXAfd1cdHkQSmp37ihVETA+bMe3qPClD3YThL/poTXJF0qGAGxViL9w5Gwv76d82EwCnKeOwrj
MgY5fWnQG4yy7krpH1ggqzZlloNdhddpYOAaTVdVPMdexaZSYvUafvYuYbwW2dLq3fdyYNKT1Io2V6H63wgKoXbT/ZVCDue/5dxF0VHH5fxnckI1i/bOzDo7hjcWHXWn
/NpjZMHdA5MRgX4htPt3vYNxF05+fMMIhjTy+zEu7XtgJM5/BmFCV37mY4767vPIXIA6IN7aK96lFqPI7XaeZoWm3kueHxLWvT6Wf6AeeRrKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiHIHLql8/FShcQ41SVHzY3bMlrA6kAKGmalSZre6myAHd8j3axqQaW8FTnWHHmHrRoTIWzPbNGKz92hyIJqibP00Yuv0O/po2woqlrVBpjas
6urTQ9h6dr/rxkDOao2lfCjBXTEgUERnGbUa0Ump+WaSNw09cGng8UC0zuarcnzVQ/kHdNL/8EuqgM3m3ww6WdsSlW1oJVb7P0LpuQJagLbWQN5NBJ63YRSJ8xjWyfzc
xfOL6yVsaWTlUXlqc8xSFUts10MoVIJgrWj0RzaQCLQ8EyhID5H/ht56af8vWeqFA5phgSXM6O6ZeT8uyPcSu0DbhtWBdAzEGqD4uoGyp3KHWZVFN1C4ZdsqpdxEhvEc
Id20p1wMJ2gcq2dHcZluQ94ER6ENG7m0FDD1bgBFTDorT0IBoL4Z0+hOhwgDG/l4R4Qk1eZA1wnmTX0SJJAkPG2aGZtJAW7/hBnchCAxhDie7j1ugJyVc2hfe6Dgaw85
OphwATLtaA5C0EoIoK1V9OF5aQkxrURn7PVlSLbtU79FTtzj4ByygKnyQoSrGrIyxCPxV7lucI2gInekLROvH+QicRefA8Lj/is1zeV0wMORpQjoF0MHhwFqQCq8NNbS
4L1dGcevcyGIUXfMoKeherFSkEQchg0CCKwa0FlvnOoSRqiVp9bf6hq6IpjBQBhWjhBUmbNndoysNgpFTCTRQ85yydRQ37QSt1uZKSxAfPeorqXdKFuVZY0h1osc8y5S
NmAhAFCQCeK4ksHy1Du0uUO+s7ZVVugJmifn0NlOoN1U6co60/5xo+OxKJHfFKodcglJfEMN51610fgkySO2xtKPFPNN4I4HIDZjoE0FIJcdcVRoF1w+oVewStREKQOM
EQNeT0ADXzgBH+YSSlEgOmt3+HddpNoLrTwrdq4Aa/x0QylWTT+JUsH9dzyAo74D8eFNKFJeoumEjSJXIZ7AiiqPZvSsJfn1fRBz/Evb+4phUqSvC6EjN+JM1BloexxE
EYUBbJ1peYPMQtNBozxHh7vXxXn/bKlRMnFeWWj9YpbS9n8LkPi7FXyEZHTrIDFzrmoqlOCgfL5bckf5a8wiBUmV3UcDeLGhA/7PNcP63UyrpY9OqzrTG3VR9UcCk3LY
nreOuqgKTuhm8gA8sOhYIZ2ZrLqi+pUKtkYfl/1vm/VAyaqwkAgzq4ApJkwTRqQM97B2JehCxg6I01SnzShy2MqIJtEmvYeBjKtfeWMCbYgzTHwCfWRG408mCWP0CV5T
WqXK86qjY60oAmI0XxW2CwpauZOF4j6D7dHbJNYiI+H9rZ9K2Q0B6dykSwyeg3DYEHR6/kXGSvgBo8E9CLDK/8qIJtEmvYeBjKtfeWMCbYhpbA9bK+Xi98MU1HdYmi9D
9s8oW7v03dmaaynex41gDvSilCo+nOHq1vw5gI9W5BGBGsicGBkPX0c32PkFnOejKqMw6NkQrfbd7jaT4gxzLMK6z9P2mIN5oMzY5t8IlwmMb/a7iO5xuloQcxWXFwIN
GbEKAdFtuztr2Ylf51jKzRsKKRvNDL73asEZwuDXkixmgmpNWLWJVEUhiZ2nvig0EB6WNsajwUj/3iVxHSq7S0CN/ND3XZvaB8pjXVLWrgOOId7m8/+E5wzNChrkA01e
84izBkWoasb4tovD++gOScC95JGGR998sMpmNeScrVOeQ8QsxJAEjcphVGeA8TFGELLu92LMd6h28f9Lmpc9wcqIJtEmvYeBjKtfeWMCbYhcFiiPOQcHvw3+00CUmC9a
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iqk0+QnuAP9cZSNfk3qrPxV75GC1/5ojCuIkaaOCknpFfERtfOPf03lhTZXmjLajDF
vkYLX/miMK4iRpo4KSekV8qIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17uv7gXKS4CLeIVJvviXVr94iTzaeBQzdz2bF8pd5cNDI4KHCGu85PX4u0hMct9+zl
iJPNp4FDN3PZsXyl3lw0MsqIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N29jmB1bs9cP81EWpN/jx3+wP81xEf/yCOtXCmcu1t9K6EyFsz2zRis/dociCaomz9
A/zXER//II61cKZy7W30rsqIJtEmvYeBjKtfeWMCbYg0WJUxO/J5Lv4jdnSpFDRf38rKnifycwHiXqkTuDoWWVszMaq6ap4QGUdSKFEVhsV0/c/CEL3KOeNd6DNdwbjh
Dk6zYFbXx6Nl2SilnyRtQGhIFomNBuUYuJtKSRJNDP7KiCbRJr2HgYyrX3ljAm2IMa256YcMC0oL7E2ZUaa1gZz0zE1BFXlYc9e+rEK4o/n7rICpy6vrQuFpgCGDT3b1
yogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh2pA1nVT/5Mu2lBFAde4OHryogm0Sa9h4GMq195YwJtiMdmmFZvPoDIoXUrUt3aIb+W6Vn/b+PuMxPrBA4imxr9
uPRkUsxt5NISJJWm6J0GUMqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqhgHU6tMXhWGtdTKOKVdJ4IMqIJtEmvYeBjKtfeWMCbYhcp165y5a5xLjxKvNjW/gD
STjFH+mb/MbkfV5ZW3hf20EmaUhTtqNXgLqditg2MJfKiCbRJr2HgYyrX3ljAm2I0vZ/C5D4uxV8hGR06yAxc0oBELkgTYRTKQljRiUfAoVcNTOtCc+GcEoyWXd2sbju
0P1z7btnOqj0MScDpSTFyjooEVAxespFc0Fkl9ViJzE6bxu0atQSJvviQoUXQqUzyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60++9ddUIVHmNFbfzkzmrck7z
p96W3VtnIC3fvWoipO87QuKStgkrZ629oZbxnB8ICv+2lI06FVws7R/e0mm0UfEWgKY3HOKtNh3t9dyzixdUhMqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
satE87EvVlmGcqF1u9dvhmwwxEkOuSmVfXhM1MA40otBHZ58I7/MXFr/Gna5HWtwkSZJhRovzXpnHHpbujOFWmLZEhaR1plDzfRfKPADeypEZcG++MHBA8xUNbXYmCNX
gRrInBgZD19HN9j5BZzno6Nqo6YHwZu75vO8OVH4V3P9T3Lp3qmLK9Ao0TJyWfuv5CJxF58DwuP+KzXN5XTAw9lCV0UafUhRzM4chONDFDCf+SWWJUsyFnlGIDK0qiq0
/JkbSQkpJ2qeb/ocfmMCUaBTe4B3k/mbHjIUfqo67SJ6y9i30K97OLHh9P33Lu8lKYzZul8zVQl9latWjvxDbo7iQ7nBaKh+iDx0aaXgHgBbzQIbnjnQSeLTnCw1O2W/
I6MZOJ+JU7iLo+xdUSBlEsJMBRG3r3K7H+sBRixxseKeQ8QsxJAEjcphVGeA8TFGAkzUKh+ZI77hc6HeH6sjhbBAgW3YHXeCcn5PVWdi1vjw7haRU2FIPEVTdfREZzeL
JKpEeE9iq+Ri+S8BxWEOuF8rOibEnWG2W0adFG01S/htolL4LqwDdXrc2Mg589fD9eAhsbYpcvuVPp86ImPIqquJfDX8tHTdjlN1M3XhQyFgve8ymNkD947ZoOaO/rwF
5fJLrZvThQEOQZCsEj40lDCgwAnkpfV+pIyXuowajgRZOqHzYc9BngUWlAynZQ9WT95ue6BORD+9cMb/oPuB2oNxF05+fMMIhjTy+zEu7XuI2yGewAgHRVNkLO+0IEC4
ULIJMn+2MkmXlNl3Vv3yFkmV3UcDeLGhA/7PNcP63UxJqsVbVLvGRAyJ2WuAecKPY+JMehL0jLBeHC9XZoz1XsqIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N2
oY26KE0z3yVq2wZ6gHZmTNN4D+wHk19YOJEoBAac+tXKiCbRJr2HgYyrX3ljAm2IkbBKJgiwwqdoMivfKpshCEyQwht14NOkUF+6aoVut9TKiCbRJr2HgYyrX3ljAm2I
0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+i+xh5LTFJRx7Fg5U3IXHtIyogm0Sa9h4GMq195YwJtiOyH3EcaH7sgrt2Mfu7haqR4cy0i35Nw7ClctH5qvnuy
LmKRiI2lIu7X97POMWrj609AHUqNPiKMXd6TmqYHnDE8EyhID5H/ht56af8vWeqF11cAtaAO9BXMvrMB9ZhZlUTogJKXOvj2i9jswBX8gR01O9BFyh+oKBE8Rum4OZBp
Rh7rZFoDrhab0P5H8Q6h+ZewoIPnpv53yku49gQU9xbeBEehDRu5tBQw9W4ARUw6K09CAaC+GdPoTocIAxv5eLYEu5VV6RvRfKX0i2y39rtffjDKjWFZ2z1UMFrVfr4K
Dkn7ihq/0iEIt6k9El9y10v/5Bu3sM5kRp3eWj5npEcnordGSFLJEKe9MCJqY81ayogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBm/F7SPlj00QfEG9vyk/p0+
8FpnaOU8oOxbgtDgG8ilO7JeLGLjyYa1obazmi9u25TpBPsLc+YXB1Nh77ougkYJqDuOw8l2Gf6yv+JRmGt4hjLOmKfN7GxIo0j1RZbbETASRqiVp9bf6hq6IpjBQBhW
1tPwbh0rHsqX28rLT+OtJ1Zqk5Dk5jsxZ+awdOF5hxIBbnrRcv02JPRKCRpsm/DQa21ojStDfqMIR5tPLKeE/w7f6diZ6LcPrbzrI1dj4T0uYpGIjaUi7tf3s84xauPr
HnxxE58x7qzsr23/eeD5yl5/vxI/XqEmevWJotB2YdfKiCbRJr2HgYyrX3ljAm2Ix2aYVm8+gMihdStS3dohv2GIERP8AIhEEaVcNxRXd0jzwkqEkSl47BHEu6PiJz9F
yogm0Sa9h4GMq195YwJtiBXSZE99vYuwjp4TNSmMSqEqdeyIf9wEYO1heD/4OzvByogm0Sa9h4GMq195YwJtiITIWzPbNGKz92hyIJqibP0C6hxlxGIQn2yBxu8tXdq2
wu10agnpq9ybSsPW9UOYxTLhxmhYqgtFWuNBznYYskvS9n8LkPi7FXyEZHTrIDFzmUDYNE0/f+Eu12vm7ePmpsqIJtEmvYeBjKtfeWMCbYjQ/XPtu2c6qPQxJwOlJMXK
ceBnFCe2zaYhEqGkcX2ypQZEG+A2CTidlB3wvHMt/bLKiCbRJr2HgYyrX3ljAm2IQMmqsJAIM6uAKSZME0akDFQRbIsS2Idlh8VsoUqqEEOn3pbdW2cgLd+9aiKk7ztC
4pK2CStnrb2hlvGcHwgK/yVuG9Op3VuX8NcJNVTabNZCDY6kpPPo85HB198p+T1VPWzu1WVz94cYTu3XYoQ+FYmvX5jRYBoyP+S0/fQvdRqpI19qwryT2npYg2oNkgZF
bDDESQ65KZV9eEzUwDjSi0Ednnwjv8xcWv8adrkda3BXVN/cAfQSP4IKxC3JwOR5yFKeMq7K5IySuH/TRkl1m4O5HR9IKDWQlW73H0bIJSJ9SChKNknSZ8s69N+tqhXO
qJyIFPds3j4XyyJESgGsqv1PcuneqYsr0CjRMnJZ+6/kInEXnwPC4/4rNc3ldMDDvYV97WOw3QgbNDtAPPiV0u8TbH0p2sD6dONfI3aiD1j9QHt/1z9lEtaQRKL2awxs
6cdV+3ONhDnp7Kb9AzvcQugJQn/Jc8KkEKndei67Hd8pjNm6XzNVCX2Vq1aO/ENujuJDucFoqH6IPHRppeAeACIEBeGptREpFM4lDaupomlIHqOfEHsLTpHSbi5HZyKy
3W0mzfqhJn+IHnJip+g2dKGOGRbTFlHiOvUQpjJMgs1CsQW5q4MhKtZrSXHYjiznsECBbdgdd4Jyfk9VZ2LW+PDuFpFTYUg8RVN19ERnN4vK3Q5jZo0ofSaGQHEG8LXk
0/0JVm027GiB5HHf3+3nce0J8Y/YkN1r8cIfZ/brhS42ZZaDXYXXaWDgGk1XVTzHK/tnmmJQZ01gcWzp5jVjvWC97zKY2QP3jtmg5o7+vAXl8kutm9OFAQ5BkKwSPjSU
JbrMmTSyj9n+Q7wjTtehWoxLBfQTrASXbWueBcmb4PBbQtbEx0pSk4+HSIGt1s3jg3EXTn58wwiGNPL7MS7te9rEnm3li2AA5V4HmErtasFQsgkyf7YySZeU2XdW/fIW
SZXdRwN4saED/s81w/rdTAqJrloSNP0zFCLM92m3MQDpihAanr3fh1KE+ukRthhFDeBYzHp6a9CkETVhD0tZu3IHLql8/FShcQ41SVHzY3bMlrA6kAKGmalSZre6myAH
03gP7AeTX1g4kSgEBpz61cqIJtEmvYeBjKtfeWMCbYjhhg2OPebVP/2RZKSiMqXL8LwxxcpN2iOFoHhbtf8hKtiMYD8eF9P3gXRMPHskkYjTIZGc9kTWzrYMDyDvnYgc
kjcNPXBp4PFAtM7mq3J81b7GHktMUlHHsWDlTchce0jKiCbRJr2HgYyrX3ljAm2ISbW4FPrgHKGV0fJhriJU1W0xohjSzRs8thLEX+w+oH+ZfnCCHqSN+ERO5Tzjs0d9
T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCDkF/pg7pGqF4RgjzHHs4KtBCSAeGAmnBJ2ZpZaneHbjpVmPRfgv4SEuX/I89VNiOI0sTxSc3Fb+JQMAdAnjo/J
vxe0j5Y9NEHxBvb8pP6dPhDJZC76kMgXde4b2XZr02DcD8dBQBgcZjBz164qcx/8/ef8LckCM5LbZZLZX6BZ9QqOyhoKxJaGCt4myMNaNZKihA48bc5x+s8XQQVeUTR2
CL0lFgs+zy6GkVajyRvIAtxNVTyrJcJJNJwB/K0ICjXI3jXGSaLMDTPJMu0+Nyg4RU7c4+AcsoCp8kKEqxqyMvxe3ys/Z7A0Akzc0zSOQD8CD+Ub2TcuiMyZVl6wfe9+
VD4QniDKrQPTtDT9FM+FaF3fzdocUbykuhHP8KYqAXWfHGHWXpSTo7z0ZoJIsD00W0LWxMdKUpOPh0iBrdbN4/rTHr1geMtXcmkU3abg3u6Z5WxADmUCAyV1dgP3rTru
yogm0Sa9h4GMq195YwJtiKpk1g1+NFLOKFDw3DyKaVTKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhZKODriqAGJStbrevKmGRQ
ho4Bk3CGftO55JtjjGCmgMqIJtEmvYeBjKtfeWMCbYhZ7N/dC6FLP0cRj8aPjc9X0iOE9Q4MxWz8hAM+uRHc1cqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
sFCxlL+i3dTIqtDlf6gD7riwuC6l8+ctLpXTO0j/XMRZDyNWIi63qHYJGUln+n5IOLYnzvzwmlP2wbbeF4bsNj71HTn14m81fQy/PIbQNkTKiCbRJr2HgYyrX3ljAm2I
2OXRUnXYWyKeeVYLciOgsqJ3SiBZNStaEB5FbOxR1/SI0HcD8Qjccgjlq2zw5msnJz/MOFTyU/ALkx+QR7tnOhUHqTdhzqoEUShXQZTAAU42JmECoLNUZHza0HpnqesK
Rp1Js5asDMFmrZkwq8nl0MqIJtEmvYeBjKtfeWMCbYjeBEehDRu5tBQw9W4ARUw6kR+DIRXv0Db8V0AYNCWTfv1udlPZLNrWsO9oIpTwPj7KiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiPwC1hyy/IvhypcOsLLeE1E4tifO/PCaU/bBtt4Xhuw2hc4jSwzDsq2W8fvr8FGgKtM7DRjPoSaQhCOO0qfyKMDiyXGgez6OzrokqSWEOhFc
yogm0Sa9h4GMq195YwJtiDvJekAVMZ9743A1UAbSS0TKiCbRJr2HgYyrX3ljAm2IFQepN2HOqgRRKFdBlMABTpzc6TfRDiWl6NCjnP/VxG8CjZHY7aFSwovqEW8xgJlw
xuZfIvjJqt+EK/mvsE+yQqpNgDYGcjvWAWStDOu3XUXrfJIOBCQYW3JlVVDYsS0UPbiZf8GzbbDB7fRbIAsY2ICjv0vYGEGhB3hfzRYrxHXKiCbRJr2HgYyrX3ljAm2I
qd80UxWhDv9pm7H3Ktx3+zi2J8788JpT9sG23heG7DaFziNLDMOyrZbx++vwUaAq5vAaQVB3pJYyK1G2e7VryXivj/guzsImM1U9g1wgqM6yew+YKKX95bc4k7nJweMK
XY8hfohMLH7MRrVnz5v3cZ+NgnnNe8IRCQy9tIWQOVwVB6k3Yc6qBFEoV0GUwAFOKaJiHMDiUQaJQgKTBOvJkQKNkdjtoVLCi+oRbzGAmXDEgsQD/dD89Tp6T1lL4YkE
1IeZfald682iylfJdWxSCd237B4p9fDB0WZsvqnbvU4ErSWsFZM42Mjk+ng2x7v7bfLza5EiNVcf9E6xuzYnAIRygZs8gC7ePWhWznkiF+RPFmmWrsuva6ex6XdAbcat
ktHrT65PHg3d1uYB0V3mfRW1HNBoz9wVrzDRu82XWYdg5RaoiTEX6pjSk7CiwTUzPfxQezN4tYR/9Kyi/Y9D6E18NiDuYCf4w9EDbaY6+W7KiCbRJr2HgYyrX3ljAm2I
F/js19G1+Zlu9G54/8tloXqSbz16ZVJjzfHOkejbX+Wp/LwAImUCLKm85fZVYqzVBK0lrBWTONjI5Pp4Nse7+yXg4J4JxhOQ6RN58jNf42QCjZHY7aFSwovqEW8xgJlw
TMoX4C6LdB47Pa8VbMIEbhCfDo9Gp3AQRT3C0sG/B7y2gvw90JwDkQw0QlmSus0KQiH0lP1T0q+aS30h6vNObJ2brV5VFrRHaBlhUIR/mWI37BSe3gTfcBcgcqvFwLaI
CZhM9Y/5TBqOD0MgtkvlLsqIJtEmvYeBjKtfeWMCbYhlMJUJzBQ58itm6vCfFp07UVhni9B/BBJ5Ohb7t/ezaYFP2uVnBSom1oMBwbttk+CCkTXC9lUQBqVqT1WoRF4V
B1GM1mcHalfl6b/NuENBRCNwngnmPbnkdFnTLTNQ01jpxJ0TMHZ63tCZWLz8JjX5YuZcZvsOgXX53zmcbrTRr8qIJtEmvYeBjKtfeWMCbYjOFk698XPU6e8XRKTct61w
IKpc7sitXnFfnME6aClAoVd35wlVjPs8vylN/12C9AQBaMQceqXbNR1s3fPXvPBpXR/oZGrTmQZTHqDmvUqVBsqIJtEmvYeBjKtfeWMCbYg4QaZAOvsVW+kk/dOYU/lf
Gtqe8iE6EqJEk/oEsvXuOeFJcMVqlH8LPHKfABir83+Qqp5P6+PAEJkWh54fVse4BoMiHPw5GySYp51IAbs4wcqIJtEmvYeBjKtfeWMCbYgz0n/7QNK11DT+RKk6bmC1
g7Ot0oLiYJdZ3ytI1KeQGezxJgUN12Wk/sEe6FG6IKan1HVV+A1MfXYmt3QZuZP+yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYgcjNMIr6UOxuen9d3bDBUp
FwZbrAYkJwYqvi5vJ2unlqNXQyAz/3DXpUKKCL8MdvxHPOOE5dFYodNr4oxaBWMRy3OdJDCzk58C2lejcZTvLsqIJtEmvYeBjKtfeWMCbYj9qdN49JXpCwK+TDd2IgVw
ZMWnhSJsCiQZp9R4CLtip2ll8qPrtXSbNaQtc+aOlqzZzK2UwFCsnK4p2KfWWmksp95uCn5vV6nZKE6Pn9/72MqIJtEmvYeBjKtfeWMCbYiQENDAdsGbFa4/ZiSR2T9l
0QgdFNRYsCLXEGiwh3dXiITB+f2g8aZbnLH0ZtiMJN/6cEdjYU1U9l78zxMh+ICtyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYi625YOqziL0DXzC6PZOwF7
vaoQQgOkf5XNyy/XRWKV6/+wiGAaK9ut0YvRaPyrXUoeY7E0HEftjj4Zd/J5OgjtQYXVdxVtr4YNkXXMwczoZcqIJtEmvYeBjKtfeWMCbYhmfZDuytXCrQ8Geix8wiQB
RP8hbDTbK8np+Qog7dqGxZkxbIMllj9J6nQD/oVUPoFqPW04tT2VRqsu/BMhMijLKD0nxU+vzPTg9akYTDlxR/PlaH+v3BzWE875q8a2MSHKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiD1SkFCVAEtdUAby9OkH/xC1/+TTc3yIOB9nmyVVknTZMg+6Yx+cE/kBgVW33wZIbpCqnk/r48AQmRaHnh9Wx7hYYGmdwBmxA4BBEut8cVUK
yogm0Sa9h4GMq195YwJtiJZS0GfYOcZrQc6u6ws0ymNeeHFHvz1V33g0ps+Ljk/BDlps86NseSF//UC+KH+djUmV3UcDeLGhA/7PNcP63UxUt2XNRoOxmqfudlCHTWRy
yogm0Sa9h4GMq195YwJtiNxFE3b+K4iHfrwGIIydTIRUPmkanLbyTCNYvwetJHaiZuGWm9IIjwOEJmMEC2T2bsMSlqqadTNMLHCnksANWMCfm3IBLLZyara6E1AhkWJ7
COqHByFykjDJdGrND4gXzcqIJtEmvYeBjKtfeWMCbYgwhhxf35n5tq5O3opeVf9q8VsGJnzdvZl2nVnDVuVPMSRcdz1x08Zr2ICbDdMAnCHKiCbRJr2HgYyrX3ljAm2I
6Wf6xSYPenzXwunwtgoenIiTzaeBQzdz2bF8pd5cNDKxMGawA3NAT+Amu5bq3hkbyogm0Sa9h4GMq195YwJtiN0pz9mKF/hVVkQ31AzIulsc2rnX8uue1oA+evZh0ISG
o/12xGv+SB8cJ/LwfjLUejDNFD8gQC7qU++CVTMiniyuWx9flS5B2tUtGZ9aRgmlxg7m+5aCTKTNvlkcTmC0eqUeIwrfQTDM3zgfMq4eOFZ7xqCUNVolHb1aY0m/p4+L
txqHizodiXsdx+fkUX40EdYNJQeGbLiXNpanKsvD6k1Jld1HA3ixoQP+zzXD+t1MjYX4XLjun2wh3SsX57xk8402nP9jzzlfQEGefwpwncjLq4qCTxktIyblMQhAmbCh
dG8cFsWcVMfy3KpdNwWSCIlAA/18cor03O4SdSpFcILxm9Gdd3B9P8Jpq57h+ON03SnP2YoX+FVWRDfUDMi6W/VGnrA1nAcyrf8gByX7JMuGlB0gAKu9uTftf9ap7WXT
jYX4XLjun2wh3SsX57xk8xmRuQulVpEVtauXqPxevylYpu5vPRSDKBBaEvE/hSoapR4jCt9BMMzfOB8yrh44VnvGoJQ1WiUdvVpjSb+nj4vCNU2BJNFSQvQSJJgsBGNm
j0SkJkrb4pVoTzDHOoaVPUmV3UcDeLGhA/7PNcP63UyNhfhcuO6fbCHdKxfnvGTzlJ3c5pwy+8Ywbc3Js4SRBdfNxhHNS7ui8eEpPYwa94cXJEi08vZ9rXqEtG9uHZD6
d5X6rN6Vxy2D3hLOMefQW0mV3UcDeLGhA/7PNcP63UzrrsCKD9x7qGx4Q4q4kDbqyogm0Sa9h4GMq195YwJtiLKHvVLnmsvoh/nPRysVIasSZs27OK/4aT2V2Ya36YtK
z5DQxMYEwENADaNiC9pvotnMrZTAUKycrinYp9ZaaSyTfZ7lr4cO5fuNEfX94qZSyogm0Sa9h4GMq195YwJtiPg3ra1WDKOP931uIhlUQHF3pqShCXHDzJd+wYBHV6dS
ctWYjJ6LNvHCWwyn5jtUtLoDZElcj2/GKFGCFZYUI/C+I5RtgdDIyt3IhpSSZKgx2IhYvXxemcZJ6GB/Rh2d4MqIJtEmvYeBjKtfeWMCbYj+4cd4u5q0WVxMxtspIbru
yogm0Sa9h4GMq195YwJtiEXfqrGTQghLSkc8wiVaALrKiCbRJr2HgYyrX3ljAm2IjDmYPt5UUsmdgOP9xwM5tji2J8788JpT9sG23heG7DYdBLynpxK/Je/G5JmdVeLH
yogm0Sa9h4GMq195YwJtiHswOCGayFX/Gmrtd4+JwwCBcW6U4hfHM8TeuEhmvHBGLnBPLbCjOLf5W48WzrdlR3AX+1zx54GE6Wpw2PFgScGt4GJHMPwvhMmbAn5+nArK
t18CgL+5iGuF8GzCXIFql4aGZSAjySL+mbE15jlpxYA9cbnMRKzjxja01XCNxxLfThieUdEnWVjxw8wapHS5hnE4u1EH3mfQBHgBNfYWtem7Z+KM0ehKa/R8Xy1wWDA8
lWyBJQMEaZO8ltp9L+Z2tQnoid8KBMDRENdJS+fpF7UCjZHY7aFSwovqEW8xgJlwWMW+Z9Yub6Exshrd8ZM7ZJ8dpKlkm5zueSmnBMeRvQCUVNyq2AQPD9kvJB4JjOsp
IV1Hafe/D/YONJfZo9gUV9u4T4ta9Vyv3W9xug0gUVP+jUZ4Dg33AmKe1yvibhKt3tg36JZIjTN8D7VQ9R/Vsl2PIX6ITCx+zEa1Z8+b93Hw3LoFsIfSx638mywsazh2
lGvRoYzHVDQoa3DsAmLyrsqIJtEmvYeBjKtfeWMCbYik3+2wZvNVc1qYjb+TDgaryogm0Sa9h4GMq195YwJtiNwjRhzctKpJwQ2CsTwsmns4tifO/PCaU/bBtt4Xhuw2
YhiRggejoYHv6vFEMznqjsqIJtEmvYeBjKtfeWMCbYivh27m08EJ94LE/av897uTKz8+1FN8OHEithDF8u+sZbrlY1lJia7hm7IoNm8ohVVPQB1KjT4ijF3ek5qmB5wx
mKF1ugDWthNttJVEQuUer8+Ak6yGH33N2+czGxUa3ktj6dpd2KYfBNR0fBwjLdqkzUgor+pCubWvNi9GR8v6xBYE9rWRMSXx5qAGUF3JGnbM1xWbAtSgUHoIcuyQ87kS
Zdli1iwbJ4xPvoL6A/SHCwd9edY91b7+iY74hScnRydMAJrDHmKVuGFnxqGbA/1pyogm0Sa9h4GMq195YwJtiOXqVA+HPfjc5jReY0a3zdfKiCbRJr2HgYyrX3ljAm2I
pNWqDhJd34Kt4/uLJYLxw8qIJtEmvYeBjKtfeWMCbYiDzhSXBFbyC/ragYHjZdZ/ooANVZv2tWFy/3q6uPLNh91daLvNXNxXiFNj+HOBmEzSI4T1DgzFbPyEAz65EdzV
31AP/06LkOpWQry2xfiRhHYzUTKn4/joLPh+0mnxIMXKiCbRJr2HgYyrX3ljAm2I4m1ZzMaTtVxmuSNJ8OjDjVCzlhBCozpTbUNadXZIp4G5dOQ7EQRA/Yb0UBPNPlvR
3MH3yNHRPOMmuAV3JC21M0wroDANtGogYx2UAaFHj/OBPi1c6vo1t52SfL66p2z6v8t1/qG2KXqIRYco6mydqdqzBEQopfOMZzDLMuMYqli3XwKAv7mIa4XwbMJcgWqX
BTRUfqB/L3hQmX5Ys0KP+fkgIJtH3AOvMfUe0OEITo3OJsXyQyz14v2Dbz0sstILSZXdRwN4saED/s81w/rdTI2F+Fy47p9sId0rF+e8ZPP7ZiEY+ifd+M6IJNpIwu7o
6Ic9+2qos/+ZkaQ+kPaXu9CunrVxnkf24yUwbNo/pBPq0KEWebp9o4S/Ms7L7TWZLnBPLbCjOLf5W48WzrdlR6HQz34W/DgROzPwAYU1Ibm3PzcpnhZ/y/C/MZicuQSQ
4UKngL+7lUHXF0NGY5e3uhYxBXikV42LmPDpp1Hkmppn0icwfq3qMmyHmOd92b1pOokRpfgaJTSmXSkVCkDA6tPmCoVQsojaaCu3y3dbGE6HzanGO4+vXTk8Jcuu+91b
yogm0Sa9h4GMq195YwJtiO1Oke9IYPfoE3oQESIhVy78VdPacW5SfaKm0cs7qAdFyogm0Sa9h4GMq195YwJtiIKlkWEh23ltQ2FucV0vNiDKiCbRJr2HgYyrX3ljAm2I
m3Yfvfg0ViQLkDJ2do3grNO669aHYhjcibvMHqfG0YV/gw3YxV0lz2HYTkiCS8MNyogm0Sa9h4GMq195YwJtiEhsI7HaH8v7mYuhwiDuLJ+EWSRaPeHN44Qhibuv56xq
Cfm8+2XzTBowM6ocCqgV0z40SZJh8I4QA/tZxC6CeMDKiCbRJr2HgYyrX3ljAm2I7k0Uwq9vV3uzLjRoyGaRn8qIJtEmvYeBjKtfeWMCbYjLXIFhKnCQJyCrZcABWo/F
yogm0Sa9h4GMq195YwJtiC9XU7ARFZG9AcHqL9aQqZ95SkuU3RHc2Ir4v+i9y/mWgmTlXh51S+UdfEX3Y/IgN26fpog5jbd3T1z+Vg/b48CBtdaRBqeOTD5UUzy+4K+A
SLXE7wNgOsZWOCqmq3y6es/gTP3kfSJxBvrcY8H9AHTbJd4h9I5IxNAMQRiKjc+3B63VtWrq06MvteDHzdIec0d+8/x0979mmloRl34z6cDrZUD1tti+UlFo3ZVlGOlZ
2uM7DW7NNVRZIe/w/89bKsqIJtEmvYeBjKtfeWMCbYjpWyZBD9s1GsVy/yZ9J3fpnNzpN9EOJaXo0KOc/9XEb9w7/5F88CKrB2TX7h7EcMZ/or96D7N8WBIZv1wdbjbF
BQHuUsgrUxgv0XDnGkF9aSYNUYo/lXQJmTOzto0jzh2bK33+Ye9chFGSYVI3XBu9qmlUgV25a/mU7ZlpoFzxba0TqLGTAdJ4F65f9v4mbqdw70Un1Q9IUc6G91GseXXA
ql1NB7U/njFU5faCQY2X14FbXHVP1ir6k0eE7v+xTir1D21LCFwJBfxr4co3Bk5li6qCfPbl59E4T9U0ypw7G3m/WNQmp0SOE6wA2gkgLvUpsBaa+693yKVXWJwNX13L
n4xSuC/NZe+K39FRp6q0k1ablOdh7CRwTzFd0cpmXPgucE8tsKM4t/lbjxbOt2VHIGjG59PvaOKsXm/4xzckXKBTe4B3k/mbHjIUfqo67SKYyBnTbhx0GYC7KDNFWIQf
SZXdRwN4saED/s81w/rdTIXOI0sMw7KtlvH76/BRoCpfv9Z3G/mipPG21j+kuDtEsL8UraaJmYyJjew+5n8HuhFkxCIZYpD/A21RrDVEI+BqeefsxlIX+AfJNXf01AzU
69zNUiOvbUD7bx1cmh+c1je1/IUWa1nMDwhA3NSNIFlyBy6pfPxUoXEONUlR82N2O5JiE7exkuxwKVV5+TkD274jlG2B0MjK3ciGlJJkqDFPX8U7Y5xSDq9ScL5Ego0J
DFI/rafonoF72qc8aKyLBk9AHUqNPiKMXd6TmqYHnDFUEcmi5QbKBriBpdcZ+ULkCcBvhCSt5lzzPQLIGQ0Epqpk1g1+NFLOKFDw3DyKaVTKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiKoGj5MN2FrbDQGGH6xddEs3c5wuSWL0U3fW+ed3JyVWg7/lw4e3tjxkHreCiucDFgP81xEf/yCOtXCmcu1t9K7KiCbRJr2HgYyrX3ljAm2I
iPRpVLEMsNUTGIZbNGHyan6tp9IGg05flg1j3Ca3fs0r30/KuFfChU2ZSxaUFP8HaKSRT0qJhCHg5+cGTpkQd4G11pEGp45MPlRTPL7gr4BItcTvA2A6xlY4KqarfLp6
C08at0eGXfiWCkpxEvgDPtsl3iH0jkjE0AxBGIqNz7cHrdW1aurToy+14MfN0h5zR37z/HT3v2aaWhGXfjPpwOtlQPW22L5SUWjdlWUY6VlnaBs0sNKWOIEZZB4ibgsa
yogm0Sa9h4GMq195YwJtiOlbJkEP2zUaxXL/Jn0nd+mc3Ok30Q4lpejQo5z/1cRv3Dv/kXzwIqsHZNfuHsRwxoMOe/1nCtA+VBdFE82e800FAe5SyCtTGC/RcOcaQX1p
Jg1Rij+VdAmZM7O2jSPOHZsrff5h71yEUZJhUjdcG72qaVSBXblr+ZTtmWmgXPFtrIrutZ+aXUanewDeNsX2I3DvRSfVD0hRzob3Uax5dcCqXU0HtT+eMVTl9oJBjZfX
gVtcdU/WKvqTR4Tu/7FOKvUPbUsIXAkF/GvhyjcGTmUMRKPyZYKcdiCuQAYuU0tBeb9Y1CanRI4TrADaCSAu9SmwFpr7r3fIpVdYnA1fXcufjFK4L81l74rf0VGnqrST
VpuU52HsJHBPMV3RymZc+C5wTy2wozi3+VuPFs63ZUfWTtyD8tuZEE+sghrlo+ZRoFN7gHeT+ZseMhR+qjrtIpjIGdNuHHQZgLsoM0VYhB9Jld1HA3ixoQP+zzXD+t1M
hc4jSwzDsq2W8fvr8FGgKmX0kTNFBR8qdN9aHdd8CiSwvxStpomZjImN7D7mfwe6EWTEIhlikP8DbVGsNUQj4Gp55+zGUhf4B8k1d/TUDNTr3M1SI69tQPtvHVyaH5zW
lGVK1XI+wt22QZWdYOOjSnIHLql8/FShcQ41SVHzY3aocSG9tWbQ+RySDvasVFRIgbXWkQanjkw+VFM8vuCvgLW0wOddxuboINlOhOxs/j/KiCbRJr2HgYyrX3ljAm2I
T0AdSo0+Ioxd3pOapgecMVQRyaLlBsoGuIGl1xn5QuQJwG+EJK3mXPM9AsgZDQSmqmTWDX40Us4oUPDcPIppVMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
qgaPkw3YWtsNAYYfrF10SzdznC5JYvRTd9b553cnJVaDv+XDh7e2PGQet4KK5wMWA/zXER//II61cKZy7W30rsqIJtEmvYeBjKtfeWMCbYjZU+BVsllaz1YDbExmovNO
ck/3YQJlIjXXC3tVn3MuAHf7h0Kk1hBXlzcjJy2iCNqYruGNFyIgiF59As7QMgjSmABL/8IMX056lYlQ3OgZNU1/dFQI+bNoTdA3CtXKYvRxHkbPKIS9iH9bielhvGtf
JMd2zGbgOY3dHTWheH5V/cqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IVOnKOtP+caPjsSiR3xSqHakDWdVP/ky7aUEUB17g4evKiCbRJr2HgYyrX3ljAm2I
S1VBvPirY4PczGpkxwLsZ5lvG1+2uzRv3xVL8IbOree49GRSzG3k0hIklabonQZQyogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBlWvb1l6ujryD5TH+WvaG71
yogm0Sa9h4GMq195YwJtiLz8tN4kGnY71INEFSPIf3AhvBPv4szoA2bQnE+kmNvEyogm0Sa9h4GMq195YwJtiE9AHUqNPiKMXd6TmqYHnDF5l4tHAQTcyKdVO4u+Yagg
MoA6GBaA9uQBG/ZusBM7io5ZNWwwJhlxgYBcgjpWTjUmllQCq/yDtYd1swvh4v9aOm8btGrUEib74kKFF0KlM8qIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N2
RPSVlqBUKpiz/b3JoD4gIHwBsaKbAXC+3OGiD5pfLhosaEUuNR74M9qcsmYa4OSaXsRYS+QJL5ncUPlXBY3+f2AMhM7uGrm8FzWxlTypAgzKiCbRJr2HgYyrX3ljAm2I
9eAhsbYpcvuVPp86ImPIqquJfDX8tHTdjlN1M3XhQyFi2RIWkdaZQ830XyjwA3sqdIiYuSfoVc2B2O5pKaAfDbvcLrfHSCF+iPZdUMaRGrSjcOUA4yoCLOZPRMdCiJfz
VMaUMndBwF+kwMksXvheRqBTe4B3k/mbHjIUfqo67SJ6y9i30K97OLHh9P33Lu8lE7rddoogtB9oG/8HLCS7p2gOaAhQA9iKo8bjTaScZBQfe2qhrPOn6JSMX7HWXpmo
Fs3oYvLqcW4AD2lYVfJ/3sqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13LsatE87EvVlmGcqF1u9dvhmmE12LHyNDpAezjzvuWTsiU8FU2jBh9GgvpJWjq92No
hQiw+pwOh6eYL5RiJAOADPNcU1RGB/yOhfm8ZosvZsXKiCbRJr2HgYyrX3ljAm2I0vZ/C5D4uxV8hGR06yAxc0oBELkgTYRTKQljRiUfAoX5OxCP1NYuK1rrReVF4LDs
cR5GzyiEvYh/W4npYbxrXz80pZvg39WM3vWhoJgxy/jFC07vO2MIYnCE1maStDvSyogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh0MYaNhJf+YmFRl0wU/BmPW
2bPoOpfcTwbFb0FbraCaiktVQbz4q2OD3MxqZMcC7Gegb5NCX0h2/ImG4tzBlm2A5c3YPwXRvIsngCSOjW8VY8qIJtEmvYeBjKtfeWMCbYhFTtzj4ByygKnyQoSrGrIy
NeKZW51MFiTQdEUcFvEAmMqIJtEmvYeBjKtfeWMCbYjnso3BxhIoHO8y8v7ESVCJkYW//v2fiN2kzX4QinWiMt33cmDSk9SKNleh+t8ICqFPQB1KjT4ijF3ek5qmB5wx
PBMoSA+R/4beemn/L1nqhTs9lik46aRXTkSFB7QtgjJJld1HA3ixoQP+zzXD+t1MmR759Q2+mrLyV2sSCel0znDvRSfVD0hRzob3Uax5dcDKiCbRJr2HgYyrX3ljAm2I
cgcuqXz8VKFxDjVJUfNjdkT0lZagVCqYs/29yaA+ICAwjxEjG2g/jVWiWEFoRrQk1qEjIi5CfD5kooeR/eVgPgQ4cBhJRmufOgIQJ4q9m0aySCYxtoq6vNPjQREaVY0u
yogm0Sa9h4GMq195YwJtiDZlloNdhddpYOAaTVdVPMeWsb+5A6B/yQCHmCiI0hqgBtmFHFCT9vXXm68NWnx9izhdXpyxKHHtP/UafKF9VbmR+Wek2pqJSOqSC51vvhM9
nxxh1l6Uk6O89GaCSLA9NJd+4MgSYTCU5FJ+KYWwOd/px1X7c42EOenspv0DO9xCO/Yj+KGk8Net4czuOrnLG3FTQ0gcvXqvk1d7T2wkurdoDmgIUAPYiqPG402knGQU
SJsxNLe1tOsgP/jr17HwC78XtI+WPTRB8Qb2/KT+nT4mAMUtgY8OtEXzRjopQgZdia9fmNFgGjI/5LT99C91GgJVw+T2SCumRmmJ3nG+ubJphNdix8jQ6QHs4877lk7I
lPBVNowYfRoL6SVo6vdjaHGgEgMQK3tqHmt8hD0eIXtZGGnCfC9fEfGGCSwdXCSfpx6joFOeblw1gjdWHYnG7KpdTQe1P54xVOX2gkGNl9dHLkFi/FVFijqlfbdHCCXX
oaXMr+7DukL/82T9ck0fwHEeRs8ohL2If1uJ6WG8a19g6fWv1HY5JtB4Sk7LkO62qpmqWKdJ9xKIn4qYuvwJbOXN2D8F0byLJ4Akjo1vFWMefHETnzHurOyvbf954PnK
bjDenkXMIX+wNrwmT/mzW01/dFQI+bNoTdA3CtXKYvRLVUG8+Ktjg9zMamTHAuxnOPsJ6yHEbueMn+7BSrjxMdZ++rNXae4XwkuDCUWtnXTKiCbRJr2HgYyrX3ljAm2I
bhPCaJgHQmhd4PWX/OFIGSa/7PY5s051BBxptKnoLvvKiCbRJr2HgYyrX3ljAm2Il3/legucnrZ8cbtgVD8LTG+vbnG+56nw8ORyEQdcDYTKiCbRJr2HgYyrX3ljAm2I
T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCBbHLxb7Zgm1MerXG1XrJQrSZXdRwN4saED/s81w/rdTBvswdLJ5/ZqRXAxSKjOiQ4hdfuETZkqZWl8saSYgF7F
VJ2A2BvfR4xp9dBchA0gXHIHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+Rx6ObMz/SF4CFSGAaCUQUcVyCXWM/+e5NkUlgBSS4HIUEOHAYSUZrnzoCECeKvZtG
N1qOuyQmPmCKB8+i2hMab5ewoIPnpv53yku49gQU9xY2ZZaDXYXXaWDgGk1XVTzHLTgM3ZNxbtEk3Lwg3a9e1HwBsaKbAXC+3OGiD5pfLhr9VTvh7XsToHerrnsSmuOe
kflnpNqaiUjqkgudb74TPcXWUY6udJaHG40TmQ6SxiJUTxQ2Dc2SQezl5vSWbXP26cdV+3ONhDnp7Kb9AzvcQgTWDMqpyw4QoCcIiVGWMvhi2RIWkdaZQ830XyjwA3sq
zhMomDTleYoxrGtA4QjnsEibMTS3tbTrID/469ex8AtkyaSMKcZMnBkSbMuyXRLm5Y/uUMW3YfiKXbg+oak3KomvX5jRYBoyP+S0/fQvdRoYUDF+8a1/ivEHZzjHIUyG
E7rddoogtB9oG/8HLCS7p5TwVTaMGH0aC+klaOr3Y2hxoBIDECt7ah5rfIQ9HiF7eTpWnkM9e9qRS+W2ldBabYapZV4sk686kX+4aMF3P7uqXU0HtT+eMVTl9oJBjZfX
lIpI3xEqp8DvE9sB13S6/GmE12LHyNDpAezjzvuWTshxHkbPKIS9iH9bielhvGtfB83g+X1b/20MWatO2nF7yVyAo07Sdyc/JLkBGj7XNPynHqOgU55uXDWCN1Ydicbs
HnxxE58x7qzsr23/eeD5ytXoAPbltQKaEHoSqp1TNi35OxCP1NYuK1rrReVF4LDsS1VBvPirY4PczGpkxwLsZzj7CeshxG7njJ/uwUq48TH+pQ5CjNOrsEiNKj34fv+M
JbHG+TrShei7Gxuz5Y94pm4TwmiYB0JoXeD1l/zhSBlkyaSMKcZMnBkSbMuyXRLm2bPoOpfcTwbFb0FbraCaiueyjcHGEigc7zLy/sRJUIkKc2cSHcXN1M4BOIfNsNYS
YL3vMpjZA/eO2aDmjv68Ba77s/BPK13KhyVRPG2xDhc8EyhID5H/ht56af8vWeqFpcBM/MYfnTjN+ZvLX+UMEUmV3UcDeLGhA/7PNcP63UwvvmNDby730bqDNdanrDVn
h4YR/lvaYqhlthjnLjGRhMqIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N2zJawOpAChpmpUma3upsgB1KTrxHtnWxBqOCkrQb60HzWoSMiLkJ8PmSih5H95WA+
BDhwGElGa586AhAnir2bRtZqncnHbxd5h9pGqiamfnOxUpBEHIYNAgisGtBZb5zqNmWWg12F12lg4BpNV1U8xy04DN2TcW7RJNy8IN2vXtQwjxEjG2g/jVWiWEFoRrQk
KMyNAvbEdOTszf2KQxnqJY8AqjeDmGbxH1RpAqsHg7e+xh5LTFJRx7Fg5U3IXHtIyogm0Sa9h4GMq195YwJtiKBTe4B3k/mbHjIUfqo67SJ3O1aJ29U730gGfgcfyug2
BtmFHFCT9vXXm68NWnx9iyhlCkXnaPRV/R/yWO4j+sKE5TJDiIvWuuFLK16afMiSIeIg8YZdnTAxePyaHru/zUy/4VG4PBZLfml+3MRz7RopsBaa+693yKVXWJwNX13L
OJjEJ1pTyNl+buNWhdklfnFTQ0gcvXqvk1d7T2wkurf2h0CgGGsAmKr1gVPQ99p+3QREnKydwuW3mkCQ0gmg7ICmNxzirTYd7fXcs4sXVITKiCbRJr2HgYyrX3ljAm2I
0vZ/C5D4uxV8hGR06yAxc43oGX2WoIcl3ICyzmqh1r5phNdix8jQ6QHs4877lk7IcPObpLWA0HeLjvACzdt0oJyWul+lrm+j7SaWdEqKSbVUhnv0Y0xKs+KegW9Sjidp
VMaUMndBwF+kwMksXvheRlTpyjrT/nGj47Eokd8Uqh0x21lGxClIQPtPprYALnYxoaXMr+7DukL/82T9ck0fwGK1bv2AmlFkoyLvq9UvW3MhGSFkulUckraU6giPzmJl
0kONxAYCq6MUmA7NzkSbTMqIJtEmvYeBjKtfeWMCbYhFTtzj4ByygKnyQoSrGrIy6aBXgRRBGD7etqBKkIZ/hcqIJtEmvYeBjKtfeWMCbYjnso3BxhIoHO8y8v7ESVCJ
b/dEUQ3+uxt2FFY1Zb2dwfPCSoSRKXjsEcS7o+InP0VPQB1KjT4ijF3ek5qmB5wxPBMoSA+R/4beemn/L1nqhdNeeQdPM1QOQwK87cyUyWFJld1HA3ixoQP+zzXD+t1M
H4Do5XbP5QRIHRZ/4BL+OTqWHbZhHWBSAK20uvLFLTNcgDog3tor3qUWo8jtdp5mcgcuqXz8VKFxDjVJUfNjdsyWsDqQAoaZqVJmt7qbIAc8WCUD8+kYVKFzlYo/uVjA
1qEjIi5CfD5kooeR/eVgPgQ4cBhJRmufOgIQJ4q9m0aTIfhfjFl7FuzgvhEBdrNfQI380Pddm9oHymNdUtauAzZlloNdhddpYOAaTVdVPMdnnprIR08r0t4RSPUEO/eX
Z7QqaYv9Ljx0/YEtH1w+RdEdGNO5EwiGKAL8PyAj0g+R+Wek2pqJSOqSC51vvhM9QNhroIdW19SnaySHtZmVmlw1M60Jz4ZwSjJZd3axuO7px1X7c42EOenspv0DO9xC
yvI2/dZ/mQt1cpRXGGNPBVNjJN6tcHSy7WNhxKUn2CJAuNQy7CdVG4fUULlTyw+kSJsxNLe1tOsgP/jr17HwCwtyMmxmq5LN2ec1++4gOKc3pcLnZ9blzPtvrakIynYD
ia9fmNFgGjI/5LT99C91Gi0R4yyVapYZL0YYT059uCIK8AiKI29mzCpW7jADuviwlPBVNowYfRoL6SVo6vdjaHGgEgMQK3tqHmt8hD0eIXvO5j5fTtzXuCyBIoCayjcn
UBThsQjmS0ur+XHUzMZ5k6pdTQe1P54xVOX2gkGNl9fEYjvMZFCsfeIQrq0rbG6j61vvnY0x5//+0jtrNmPWHnEeRs8ohL2If1uJ6WG8a18HzeD5fVv/bQxZq07acXvJ
WSqk9BNcixaZ3y6e7wbjqytygoBgT92SUC0K1xHsm9oefHETnzHurOyvbf954PnKQcd3UT3QBs4l6MpYEp9DwnlKRnv87KxhwcJZmKMxBt5LVUG8+Ktjg9zMamTHAuxn
Lwu/LjWb9WfGDMBpEgZWXSOjGTifiVO4i6PsXVEgZRLCTAURt69yux/rAUYscbHibhPCaJgHQmhd4PWX/OFIGQtyMmxmq5LN2ec1++4gOKem+P2hFnlNfeU1FTB26vAA
57KNwcYSKBzvMvL+xElQiW/3RFEN/rsbdhRWNWW9ncEs/5+QaTWo5sL8wdEAA7FbxKYi10gIfHbaCzWpb5QUZTwTKEgPkf+G3npp/y9Z6oXO5j5fTtzXuCyBIoCayjcn
dzSZF02WNAGb1Sy/+DwWUhvswdLJ5/ZqRXAxSKjOiQ5tzoGBisywLG4NZ1GvFxZ73ZxRf6QF3YOhXQCMrdR0vXIHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+R
WeLBq0TFVdynnaWQLfUQIcHasrD7g/DN+k3AP20kBcEH+NW1NjHrI5s9sTqw6elF3YG18IQOHZAN8p80vOUtqYtga29j9WzWHanK0tEH3sT14CGxtily+5U+nzoiY8iq
Z56ayEdPK9LeEUj1BDv3l9N4D+wHk19YOJEoBAac+tV22VUlfsivRAvU1ggOKQYqkflnpNqaiUjqkgudb74TPcOcIKWMF9/YBEATAqWlQaDYjGA/HhfT94F0TDx7JJGI
6cdV+3ONhDnp7Kb9AzvcQrHVG6lC6KHv2wjgRL0b61pU44XP7LbQ0qpM+SrH2CV43dghmcK1x9mAo5MAj5zqzIICtUaXATIf11KzYbAa4521eG+st2aSJ/MQWKbgTl+/
yogm0Sa9h4GMq195YwJtiCmwFpr7r3fIpVdYnA1fXcvjL+h7LZSvywpBwFYS37CCOm8btGrUEib74kKFF0KlMyrwJ30n5KU677EG5Q/JndwEdB4SCYWlTZXahmtbyiu0
V1oe5Eu5r/e1l98li149BTPq2U9Gox8+7IsXEKhlBwPS9n8LkPi7FXyEZHTrIDFzwyMuJLwZCciPSfV9y6IaeWAMhM7uGrm8FzWxlTypAgysD+Mswa+YZU19VKqRMUbv
H+SKzx728+3vqrjqrX+uNmYs1XNv7ANxadjjWhu08mlffjDKjWFZ2z1UMFrVfr4KVOnKOtP+caPjsSiR3xSqHS/r/Vx2xS7f8cXo2mKf6rl5SkZ7/OysYcHCWZijMQbe
ncBbaCvUZbZ0R3BeM75ZSltdDv0yE3byUoH/sNuz/KfXT4ohewVhM4bpvRq63Zq3SuRgEPcZNWUXRsTWxU3aGUVO3OPgHLKAqfJChKsasjLnOlW9iV9ThBryCz8N8tWB
2bPoOpfcTwbFb0FbraCailDHbpfe1euVF6ljsJs4EeK+3/HOMBCyzHRWLdfnEbTcZS9eKDWGJfKEOP3iwhVm+OzbdcXOoLVpFJpizwq/ihN5l4tHAQTcyKdVO4u+Yagg
Ku2SR+o7BbKGc9bqEtixEEmV3UcDeLGhA/7PNcP63Uwb7MHSyef2akVwMUiozokOXItzf0GDP1CzUuJYqmK7Ct33cmDSk9SKNleh+t8ICqFyBy6pfPxUoXEONUlR82N2
BgFkoZbbTLQ27IEut7gPkWPxMp6z+LceZu6O2FcwjhPw7haRU2FIPEVTdfREZzeLn8l5SSf48TKc4bTmBS74BcryyhxHS/ja4e5Y6XTAw2nKiCbRJr2HgYyrX3ljAm2I
9eAhsbYpcvuVPp86ImPIqnsSE49SeOxuUr4WqadkYOYGRBvgNgk4nZQd8LxzLf2ydtlVJX7Ir0QL1NYIDikGKpH5Z6TamolI6pILnW++Ez3ET8fXZPNKFOVc1yEto+NN
yogm0Sa9h4GMq195YwJtiOnHVftzjYQ56eym/QM73ELXrd7RvZyz0ef3vEOF9GOoyZE8d/Myari4nkWYlJSDYUC41DLsJ1Ubh9RQuVPLD6RImzE0t7W06yA/+OvXsfAL
kEhE+JscsAzzIEdqIdzL7pd+4MgSYTCU5FJ+KYWwOd+Jr1+Y0WAaMj/ktP30L3Ua6f3V/kQEY/6qrDOKexHP33FTQ0gcvXqvk1d7T2wkureU8FU2jBh9GgvpJWjq92No
caASAxAre2oea3yEPR4he0L0gP8gcvMpiCB+jNz/IZsmAMUtgY8OtEXzRjopQgZdql1NB7U/njFU5faCQY2X10LbEX5u7FS0vhDyiIJuBn1sMMRJDrkplX14TNTAONKL
cR5GzyiEvYh/W4npYbxrXwfN4Pl9W/9tDFmrTtpxe8m6msi3Hk7IOPKuRP3VV3B/g7kdH0goNZCVbvcfRsglIh58cROfMe6s7K9t/3ng+crl4X1vXI8Z7zQaveu0jV4Q
lZI1zb/3WoHNywl6uq4IuEtVQbz4q2OD3MxqZMcC7GcLMuZ41PVTfWlCkYl4FVp3/e9qPv5HYAN+nGJsjshrtaY5XJYGnz77Iey3via1wNxuE8JomAdCaF3g9Zf84UgZ
kEhE+JscsAzzIEdqIdzL7uTRVL70LdkDJfOfXIYV3ovnso3BxhIoHO8y8v7ESVCJpWIi+u5mVmkEPlm84lRPss4fYUcLb/frJv7cbFolrKm5FYt8YrWlgrxPqP1u81KP
PBMoSA+R/4beemn/L1nqhUL0gP8gcvMpiCB+jNz/IZuRYoq8f2pPFh8H+ZTpStd2G+zB0snn9mpFcDFIqM6JDlyLc39Bgz9Qs1LiWKpiuworZxlArG8334mvAHkdgBU7
HBBXVMwMHzBKhdVnmXJsXwYBZKGW20y0NuyBLre4D5H/n2cIfuPMFsacKjOBei8K/3Oi1Ls4Vq0ZvuMlAYeTiwQ4cBhJRmufOgIQJ4q9m0Y8ufM3xLbfNq960wSkVpTV
xlixEaAG3kWLAToVwmaNGzZlloNdhddpYOAaTVdVPMd7EhOPUnjsblK+FqmnZGDmSJhpOFU3JEBDrxHqs9QEr+QicRefA8Lj/is1zeV0wMOPAKo3g5hm8R9UaQKrB4O3
DeBYzHp6a9CkETVhD0tZu8qIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0iokBYold5l/ZqxU8+wmRxbwJ5mUCE9S/oWA/UXCK8U5doDmgIUAPYiqPG402knGQU
SJsxNLe1tOsgP/jr17HwC52JdMGWhfDiEFkH1y3BaFfKiCbRJr2HgYyrX3ljAm2Iia9fmNFgGjI/5LT99C91GlZytaG1yVOzF/Gs9SZTbEFUnYDYG99HjGn10FyEDSBc
XKdeucuWucS48SrzY1v4A90ERJysncLlt5pAkNIJoOzXJ4ps8BDtBhJsiekfumSSyogm0Sa9h4GMq195YwJtiNL2fwuQ+LsVfIRkdOsgMXNL0qPfvLuLpw3E7fNczYFl
l7Cgg+em/nfKS7j2BBT3FjGtuemHDAtKC+xNmVGmtYGclrpfpa5vo+0mlnRKikm1yhv2DAx6htG2rwiEmWl+ZcqIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKod
w6EV46eQc9XVP+HwFSYcFVRPFDYNzZJB7OXm9JZtc/afio/cyQZh8J8K+G/mzUF6IRkhZLpVHJK2lOoIj85iZafelt1bZyAt371qIqTvO0LKiCbRJr2HgYyrX3ljAm2I
RU7c4+AcsoCp8kKEqxqyMtJ24oDqv4k6s5MJkTOLPZzk0VS+9C3ZAyXzn1yGFd6LuU1/Fkfj8626MFP2QYstQ8MOQGkwwy4LdoTLFAv+4kCCAe9FCVw54ZhuZT1+mcPj
T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCCIrxaN7MSSucvhOpbCqrGPdzSZF02WNAGb1Sy/+DwWUqoTeKc3MfpwxlYlT8b2xwxXWh7kS7mv97WX3yWLXj0F
VmqTkOTmOzFn5rB04XmHEnIHLql8/FShcQ41SVHzY3bMlrA6kAKGmalSZre6myAHykroj/7y3vvWkFuynJIk79ahIyIuQnw+ZKKHkf3lYD4EOHAYSUZrnzoCECeKvZtG
RjDG+XokHEhjKyrHdAQaFlMaEHlsnQsQyKZVFILUEq82ZZaDXYXXaWDgGk1XVTzHit9xbuRzVRIvAqg20vaBds6JHXwFipV4yRzFi7B2sqENa53XojgZwereuGg0aVM5
jwCqN4OYZvEfVGkCqweDt6WRnKhK+FRF8UcAIoQlSvDKiCbRJr2HgYyrX3ljAm2IoFN7gHeT+ZseMhR+qjrtIta+KD7V6s6eEW+LLtrtVjghvBPv4szoA2bQnE+kmNvE
aA5oCFAD2IqjxuNNpJxkFEibMTS3tbTrID/469ex8At9XYEn6+8omyA/fG7Y2d+3yogm0Sa9h4GMq195YwJtiImvX5jRYBoyP+S0/fQvdRqaFZe5a45cYyMO1fY/SV15
Om8btGrUEib74kKFF0KlM5TwVTaMGH0aC+klaOr3Y2hxoBIDECt7ah5rfIQ9HiF7j7Ls7HsreVSa5HrOSLzm/nJjQqQZ41m7EFvfmrlGJQGqXU0HtT+eMVTl9oJBjZfX
DbiOsiURLiPQ9Ixom59nmmAMhM7uGrm8FzWxlTypAgxxHkbPKIS9iH9bielhvGtfB83g+X1b/20MWatO2nF7ybaX9Q0whM2f+ji9DSdAQs4EJIB4YCacEnZmllqd4duO
HnxxE58x7qzsr23/eeD5yv/UNOO8kR5pHC2se/HweejIx0wA3aysTt8c67nPN0YsS1VBvPirY4PczGpkxwLsZ8iXy6HPPTxxwT7eqx9Y+3+Kq59VLpM5SEI2mM4luCdO
30DJYRfZv9E2xOEFlkuz9W4TwmiYB0JoXeD1l/zhSBl6vAbZAiZwKMo09dnN6/XLJXb1tVaGMvCbYBvv6uo+TueyjcHGEigc7zLy/sRJUImjbf4MF/0/CXFqlQRluXZW
4oya9w9tWvW4KHP8ZKPv8tP0jFjtFg2uK6V6Yc+P4/E8EyhID5H/ht56af8vWeqFj7Ls7HsreVSa5HrOSLzm/n5VqGEGHlrdJ2LITx1lDH8b7MHSyef2akVwMUiozokO
iT+WiZxsKDzs0UTeQIN/Sqg7jsPJdhn+sr/iUZhreIa+8Kowfz55NhVL3/yHRf5wBgFkoZbbTLQ27IEut7gPkVSpDryXTMXbfvbxU58hF/U9i1mOwA082XBJ/EeklfyE
BDhwGElGa586AhAnir2bRsX5LO+EbzFjMoZKbUlUm4Q1DsJRphpuLLvoXLAo1B2sNmWWg12F12lg4BpNV1U8x4rfcW7kc1USLwKoNtL2gXagb5NCX0h2/ImG4tzBlm2A
44cSrUlay67VwDQg5SUqRJH5Z6TamolI6pILnW++Ez2VauvW8EUksWHn7fVArnw3oaXMr+7DukL/82T9ck0fwOnHVftzjYQ56eym/QM73EKq2NDr8g71jrvr9J0h+pqT
0VikqnORF/odG3e8DazIZ4Gr7iVPMbDCuyMWtn9HGG+E5TJDiIvWuuFLK16afMiSULIJMn+2MkmXlNl3Vv3yFsqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
wyr6pfFQIJl8Bnay56eKrXDvRSfVD0hRzob3Uax5dcCU8FU2jBh9GgvpJWjq92NocaASAxAre2oea3yEPR4hezAMms4OF75FqRIUutWOzkLKiCbRJr2HgYyrX3ljAm2I
ql1NB7U/njFU5faCQY2X18WY87dWQw8TuAVvLwe/s8JAjfzQ912b2gfKY11S1q4DeNHW4grv3qDmoS3a/SyIHHj4XWivj1UoQxE9aC727o1BJmlIU7ajV4C6nYrYNjCX
yogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh3s8gGqpvrdfT5BNdz9LXHOXDUzrQnPhnBKMll3drG47qP2ZzmetUj/j0XoBIrVFFchGSFkulUckraU6giPzmJl
PW8nmRS1gc+TIjnbkupKBcqIJtEmvYeBjKtfeWMCbYhFTtzj4ByygKnyQoSrGrIyjvok4JJ5jxtdTRVxCygQtTelwudn1uXM+2+tqQjKdgPiSKYFKteVW/rbcRZX2hEI
ww5AaTDDLgt2hMsUC/7iQDSXFZ5fJwtpSZ2s2O47T9lPQB1KjT4ijF3ek5qmB5wxeZeLRwEE3MinVTuLvmGoINy9E5QHwrFkTmkNIyty6nh+VahhBh5a3SdiyE8dZQx/
ittRvGrXOwvDNAqnrwf5KVdaHuRLua/3tZffJYtePQUBOlMYr4/5DVlh1mkSMGibcgcuqXz8VKFxDjVJUfNjdsyWsDqQAoaZqVJmt7qbIAcAHPtJ1zzqa4OFFWvsTa3k
lFgaIwhs+0zH3ft/oKZbSwpROrCYRQK942scO9HpqGJmLNVzb+wDcWnY41obtPJpbZq+2OTrgHGsUp66ydkjE/XgIbG2KXL7lT6fOiJjyKo2vfGCRZOP5rTCn5w6+LdE
yogm0Sa9h4GMq195YwJtiGQ1KsAXKBvZU41BeqXbB0sGgyIc/DkbJJinnUgBuzjByogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0i
htAcn4WHa060ztPU1McMui5ikYiNpSLu1/ezzjFq4+uGdKOXf+3D4eGl0vIMriwVMM0UPyBALupT74JVMyKeLMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
fXwI1US6C8zsPgh8VL6iqwINWDfIV686hgH4YX/aMz9JlPaAy5vbuXVbLZfEaPG87RD/tI5p8UnfK6FXulpmPiQip8rjkGSvurHhiGgF+rDd93Jg0pPUijZXofrfCAqh
nL3Xxob8YIaf7qCcL0UNXjj7CeshxG7njJ/uwUq48THWfvqzV2nuF8JLgwlFrZ109eAhsbYpcvuVPp86ImPIqsF7PUuNTNqH5W+nRBAdPprOiR18BYqVeMkcxYuwdrKh
w/ErwKdTIBSNl/7kpInsvoCtrRvQiix+8+hfsyuorTrK8socR0v42uHuWOl0wMNpT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oVKl70i01G08GK0Xe+CFv83
axxVFBu41KnXt4hckjkLT0JyrLHFpIOVKPUMiHaY5/ORQosIdSLqoEdKclgTMH5yyogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh2kMCLGA92GaT9abq1HfC2s
VE8UNg3NkkHs5eb0lm1z9mNSjch0YORWo84SPGRyiwohdfuETZkqZWl8saSYgF7FcVNDSBy9eq+TV3tPbCS6tymwFpr7r3fIpVdYnA1fXcskIqfK45Bkr7qx4YhoBfqw
CvAIiiNvZswqVu4wA7r4sJy918aG/GCGn+6gnC9FDV44+wnrIcRu54yf7sFKuPExiqufVS6TOUhCNpjOJbgnTjGyWAI9zJW68/9P7PUFRdTBez1LjUzah+Vvp0QQHT6a
/e9qPv5HYAN+nGJsjshrtYtzeXyP962ZdA6aHsfw2R5a7ygTM7U6S9uBjpKmE2XqeTpWnkM9e9qRS+W2ldBabSZbKqDMkulM8SsRZcLRcjZ5l4tHAQTcyKdVO4u+Yagg
D8Lt/ykt2+ata7FGEh1AbdNTivR2U3mt6OblZdMp+tlCcqyxxaSDlSj1DIh2mOfzxdZRjq50locbjROZDpLGIgRbNxbxf+z96yrCQzSamr9U6co60/5xo+OxKJHfFKod
pDAixgPdhmk/Wm6tR3wtrPk7EI/U1i4rWutF5UXgsOxjUo3IdGDkVqPOEjxkcosKIXX7hE2ZKmVpfLGkmIBexStnGUCsbzffia8AeR2AFTtRJTT6I5RP35NSeu3FW+5F
JCKnyuOQZK+6seGIaAX6sN2cUX+kBd2DoV0AjK3UdL2cvdfGhvxghp/uoJwvRQ1eOPsJ6yHEbueMn+7BSrjxMaBvk0JfSHb8iYbi3MGWbYBSFuxaFpP+GH+KdjkvZkr3
wXs9S41M2oflb6dEEB0+mkiYaThVNyRAQ68R6rPUBK/D8SvAp1MgFI2X/uSkiey+gK2tG9CKLH7z6F+zK6itOgZB9kj9tJGw6bv01mwV/YJPQB1KjT4ijF3ek5qmB5wx
PBMoSA+R/4beemn/L1nqhZdfz5kSwRtuYoIjJuSW8F9rHFUUG7jUqde3iFySOQtPQnKsscWkg5Uo9QyIdpjn82ph+yUFIoWx2AjYruCXZcLYjGA/HhfT94F0TDx7JJGI
VOnKOtP+caPjsSiR3xSqHT3zOe2UCdfq4w3/9I1qGorKiCbRJr2HgYyrX3ljAm2I6hUZ8dnGfP7z4uv3Aa5g33j4XWivj1UoQxE9aC727o1BJmlIU7ajV4C6nYrYNjCX
ia9fmNFgGjI/5LT99C91Gp6tFhKLAQFqkrN6RqgFI5txU0NIHL16r5NXe09sJLq3mBnF4xSwyQWXckUvObhRgXmaq/gwnp4oQA+aXsaK7lLkpVdz/Ck7J6WDrBsWrf12
VtJrrb7moyW9w9iOzj6OU8F7PUuNTNqH5W+nRBAdPpoD/WxJpu6bRrn4hDsIxZNKsV+rFfX4G7YeBVaFSXn61ICtrRvQiix+8+hfsyuorTpmLNVzb+wDcWnY41obtPJp
zkvrbnGkwIH/ZlsnEP9KwjwTKEgPkf+G3npp/y9Z6oWVjwyx4rk7hBA3iByP1ZoCqB2l1pN+76Ef3ecKRj6JOBsgGucsw3WPoDYg3UN4RHzDDkBpMMMuC3aEyxQL/uJA
071Ryi+qiA0Hhdug1eNnNh58cROfMe6s7K9t/3ng+cpeEQpzd29+Xa185AoM5C6/TX90VAj5s2hN0DcK1cpi9B2eyDIIbmzmn2GoCA+S28QhdfuETZkqZWl8saSYgF7F
3fdyYNKT1Io2V6H63wgKoSmwFpr7r3fIpVdYnA1fXcufhBASUJd+TRMiwQq51Y/1cO9FJ9UPSFHOhvdRrHl1wJgZxeMUsMkFl3JFLzm4UYE4QpiaFgIP9Eq3NYptyVve
fWbAPcIRi1cDgZntbAj80DZlloNdhddpYOAaTVdVPMfWLi4gYaKDTvuQkrHx/FbeBkQb4DYJOJ2UHfC8cy39sri1Jd3rEY3dnrm7y4yG0Opa7ygTM7U6S9uBjpKmE2Xq
Wxy8W+2YJtTHq1xtV6yUK09AHUqNPiKMXd6TmqYHnDF5l4tHAQTcyKdVO4u+Yagg9qYieiWhKFE4U3nYKXqBiQAjbFzLYqsvIy6Fe16A/PqYd7nb05OOml55ZjGMO6Xp
xdZRjq50locbjROZDpLGIlRPFDYNzZJB7OXm9JZtc/ZU6co60/5xo+OxKJHfFKod4SKqLcVa/6YMb8cFhEBZx8jHTADdrKxO3xzruc83RiwdnsgyCG5s5p9hqAgPktvE
IXX7hE2ZKmVpfLGkmIBexQrwCIojb2bMKlbuMAO6+LCIUGmZRVAaR1raEqEPN5oTn4QQElCXfk0TIsEKudWP9RO63XaKILQfaBv/Bywku6f19eswn9HLHt1MO1f6Mv3v
OPsJ6yHEbueMn+7BSrjxMf3vaj7+R2ADfpxibI7Ia7UFzoSYDWYXE7usj9q9mivG1i4uIGGig077kJKx8fxW3iOjGTifiVO4i6PsXVEgZRLe5veDAFLNT17gcHdUkccC
H47irZgS+EA2nm7u4cefZMqIJtEmvYeBjKtfeWMCbYhPQB1KjT4ijF3ek5qmB5wxeZeLRwEE3MinVTuLvmGoIPamInoloShROFN52Cl6gYkPVz/BSVH8VlWJqQoBQAqz
NmrS0Hd6fh9XWBd76q+OocqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IVOnKOtP+caPjsSiR3xSqHeEiqi3FWv+mDG/HBYRAWcehpcyv7sO6Qv/zZP1yTR/A
AZ6gsLQS2hUt/KdN2phLJsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IKbAWmvuvd8ilV1icDV9dy0d4h67ejWrKLPf6CN+uAljd93Jg0pPUijZXofrfCAqh
mBnF4xSwyQWXckUvObhRgd8ZjqI9fp5ckCxFdC/5+3pQsgkyf7YySZeU2XdW/fIWNmWWg12F12lg4BpNV1U8x9YuLiBhooNO+5CSsfH8Vt7TeA/sB5NfWDiRKAQGnPrV
uLUl3esRjd2eubvLjIbQ6lrvKBMztTpL24GOkqYTZernnnTzaHrQQr2Uelelyx6zT0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCD/ToaQ4xdaRnVGHt84+0hJ
yQqH4PcrdglI3zOmRLulPhsgGucsw3WPoDYg3UN4RHwAhWIPaGcjKAWEO15wZvqRyogm0Sa9h4GMq195YwJtiB58cROfMe6s7K9t/3ng+cqjAEFJs66v1YE0iW6ZjDj5
VE8UNg3NkkHs5eb0lm1z9uoVGfHZxnz+8+Lr9wGuYN9dC0aaysoKaMFEtJByIXcTJ6K3RkhSyRCnvTAiamPNWomvX5jRYBoyP+S0/fQvdRpHeIeu3o1qyiz3+gjfrgJY
KYzZul8zVQl9latWjvxDbpgZxeMUsMkFl3JFLzm4UYHfGY6iPX6eXJAsRXQv+ft6yOZWpuFL37KAKDjFKRlIlHIQp5htQP28XeP4dZltkmLWLi4gYaKDTvuQkrHx/Fbe
qpmqWKdJ9xKIn4qYuvwJbCqM4sl/zqvBSvoBG8/ZT1OAra0b0IosfvPoX7MrqK067AbP7eE0lAGt/Kx24bYi6wsXJZLOX5CYy2vOpGBB4dk8EyhID5H/ht56af8vWeqF
R8M0Wz797RkQquWqd+oRNckKh+D3K3YJSN8zpkS7pT4bIBrnLMN1j6A2IN1DeER8dcOO3JTw3Qxc4GmGihpWJcqIJtEmvYeBjKtfeWMCbYgefHETnzHurOyvbf954PnK
r0wspaWVKLyiOIYgHG0EssqIJtEmvYeBjKtfeWMCbYhn6fl+GFoDhomqgm1X2FAWfWbAPcIRi1cDgZntbAj80MqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
gquHKtNqOudcluBsvWC1uECN/ND3XZvaB8pjXVLWrgOYGcXjFLDJBZdyRS85uFGB/S523EfxxwlUZm1s5z6QXtcnimzwEO0GEmyJ6R+6ZJI2ZZaDXYXXaWDgGk1XVTzH
K/tnmmJQZ01gcWzp5jVjvcmRPHfzMmq4uJ5FmJSUg2FWa1YKRXZWABDCFlnRYATyo+uvIiY/GYnLA/pR5+bWlLKst4M30vwG+y0rte+9cW8YsBNXhsW3XY6PO+na428K
PBMoSA+R/4beemn/L1nqhTiHLpNJJ+5h7Wh6lS10NLybkLKVKTSThjr6eOLne9wEGyAa5yzDdY+gNiDdQ3hEfNP9CVZtNuxogeRx39/t53HC8k90SngXIPuXw2mGsBfE
HnxxE58x7qzsr23/eeD5ypjQ0tiuNAp9szp9dU/l8SXLxKHBtsvT1ljtQATxvRZK6hUZ8dnGfP7z4uv3Aa5g3097jmH/NZ3VWrcypbH8BXmQg+6gIQByB0NisUB8a0Gn
FWxZIKJPo3U8FJciUCLQlakjX2rCvJPaeliDag2SBkXrW++djTHn//7SO2s2Y9YemBnF4xSwyQWXckUvObhRgf0udtxH8ccJVGZtbOc+kF4qcgwH0px9kdX5aYCIw4ZB
LPuy59Ej/2r8abYP90veFCv7Z5piUGdNYHFs6eY1Y73hsgeBRaLW5blz0nv6+daow/ErwKdTIBSNl/7kpInsvqPrryImPxmJywP6Uefm1pTRS6GUDc8782Nxr9qGJbkV
KeDk1zr4lzExzNvQdS6hhTwTKEgPkf+G3npp/y9Z6oXFB9jfMdooCS3fA3BDo7S+K4DvPLV0G7inilOclzZykRsgGucsw3WPoDYg3UN4RHzT/QlWbTbsaIHkcd/f7edx
I8XZSVq+8r3SwyDHpQhuOh58cROfMe6s7K9t/3ng+cqY0NLYrjQKfbM6fXVP5fEl2bPoOpfcTwbFb0FbraCaiuoVGfHZxnz+8+Lr9wGuYN9Pe45h/zWd1Vq3MqWx/AV5
0kONxAYCq6MUmA7NzkSbTImvX5jRYBoyP+S0/fQvdRpiN+39MkT/hQ3wz6nxv6vaUxoQeWydCxDIplUUgtQSr5gZxeMUsMkFl3JFLzm4UYGdDpHJrHaw/D3WdaWn9WZ3
yogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKqAH2qx/B5L2yWvUt7x/JZaAnmZQIT1L+hYD9RcIrxTl8PxK8CnUyAUjZf+5KSJ7L6j668iJj8ZicsD+lHn5taU
l0mjURa8u6sIGUa7IOUHDU9AHUqNPiKMXd6TmqYHnDE8EyhID5H/ht56af8vWeqFUh71AnViUrEaICA9w7ckF8kKh+D3K3YJSN8zpkS7pT4VBpC0h3qqEZlpZ+Q9p7Gq
QSZpSFO2o1eAup2K2DYwl8qIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKoduelAITd27+eTX80priqeGpd+4MgSYTCU5FJ+KYWwOd/FowoSf9x/Nmg8NvRekUGj
IeIg8YZdnTAxePyaHru/zUy/4VG4PBZLfml+3MRz7RopsBaa+693yKVXWJwNX13L2kFFbNZri1cSG4AU5NQQjmAMhM7uGrm8FzWxlTypAgyYGcXjFLDJBZdyRS85uFGB
3tXzwJLvbs/RgXbC/05Oi19+MMqNYVnbPVQwWtV+vgr14CGxtily+5U+nzoiY8iqgB9qsfweS9slr1Le8fyWWnztZ8/w1UxPq3rwUrUlxDvD8SvAp1MgFI2X/uSkiey+
DfQWYX0OSN0oXCmpj71l+4IB70UJXDnhmG5lPX6Zw+NPQB1KjT4ijF3ek5qmB5wxeZeLRwEE3MinVTuLvmGoIKFJO0DeYoPlDiZS9Yorsq33IxhnhUI8BgA/EhmoubdK
BAC1pKIu1F1UZ7yGeosT1waMrZyQJZIQFGiR71ov40bKiCbRJr2HgYyrX3ljAm2IhHN5hH9F82XlRyJS8p4fpUwAmsMeYpW4YWfGoZsD/WnKiCbRJr2HgYyrX3ljAm2I
LtQTCSOcbFir4MPu+NMuRsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IKbAWmvuvd8ilV1icDV9dy33PMq9hy+zB1FrRGSzVm/3KiCbRJr2HgYyrX3ljAm2I
Wezf3QuhSz9HEY/Gj43PV9IjhPUODMVs/IQDPrkR3NXKiCbRJr2HgYyrX3ljAm2IlBxUlY3dWAR6irMTNsgW0d59b5gaPOBIGTWHligEomCDMBuUX7oZMimsvwVZS+Vq
9UFXdXTkLhJvEk3v4coDLUwAmsMeYpW4YWfGoZsD/Wn7GF3hkVzKZAoM5pJGg1Hvb2VfhtZJlI+E9ouFIBY63EGXpZXyFfkhDGEWD774oi96ijmp7TPsHk8rdG838NL6
811uYMlebsgGkXlrk4FYTwP81xEf/yCOtXCmcu1t9K7CVgrO20ig/fgYhpa4+LQvxow7L245t380dzokhp4d8PZqXXjEN1yUo5XTLfRk20wEvqeC0Lqop0wJO+HpAYOe
06X8Ean2hFN0HUzx5gc2EUzVykuBbZ0/Y5XdzEZrlmdCDY6kpPPo85HB198p+T1VbJGjV6Q38mha8b8zL1whvq2QFTCYbbaJtrQ5ejLdJ004hy6TSSfuYe1oepUtdDS8
QYoAER3mW0268BpBTjkGoJcYQURHT00uizYO1XhCtaRoDmgIUAPYiqPG402knGQUGppd/bk1b+rV99JUv7QLvyOjGTifiVO4i6PsXVEgZRIc6oRLjBtWKmJpW/MpUSNh
3BYAA3Nu0BMXtZ60286uGnEeRs8ohL2If1uJ6WG8a1/7Z7wkD6b0je9oH0PHbc3FCvAIiiNvZswqVu4wA7r4sAt9BEnTleJcJb8nHeuywnY1fRsFpz6/8D42bVLsGzmh
PCYH0KIMI0Z1LAAaPDsEKGaPvrFLXr69fkq2crdPifARSMKckKtt+3ALODEHSrraxcGUgx3m8a6hR/tKenIXKO0Q/7SOafFJ3yuhV7paZj4kIqfK45Bkr7qx4YhoBfqw
3fdyYNKT1Io2V6H63wgKoWgOaAhQA9iKo8bjTaScZBRImzE0t7W06yA/+OvXsfAL6aBXgRRBGD7etqBKkIZ/hcqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOej
CaHOtUnJqSovpxwkgN5W+FyAOiDe2ivepRajyO12nmYUjclJOVXme/kqm1ln3NyiiePltBa+MRI7/E/80opPeOnPro0lhNK24jVItY11guzYjGA/HhfT94F0TDx7JJGI
6cdV+3ONhDnp7Kb9AzvcQt7TLRmxdYRpn9b++ETtzI8hvBPv4szoA2bQnE+kmNvEdtlVJX7Ir0QL1NYIDikGKpH5Z6TamolI6pILnW++Ez2jL6v4i2H5XjZdHebC+tYs
yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUZC78hPCHOnebdjSN7gozVdlwGTxSZbB/uvgmakt4kn0cH1U+PRVPXFXqvGNMvMja7Q/sOUNcTkGa/HJWED3bdx
AGIxpICnrllV6QtccNZHgz1vJ5kUtYHPkyI525LqSgX14CGxtily+5U+nzoiY8iqwXs9S41M2oflb6dEEB0+mnwBsaKbAXC+3OGiD5pfLhosaEUuNR74M9qcsmYa4OSa
BDhwGElGa586AhAnir2bRlASwzYi7xTH6Xx8UEPUKYRgDITO7hq5vBc1sZU8qQIMg3EXTn58wwiGNPL7MS7te69wR8XRHT7J62LANx09hPBLbYTiCDt8iUfqA2gWgnQy
TX0JhC9K0uU9wAlE9X6enH/OwSINmVLEOojT14nhxyTKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiHIHLql8/FShcQ41SVHzY3ZE9JWWoFQqmLP9vcmgPiAg
IAKDWCFOwDcDiXTtFLd0lTtknEBgd55k1EpaPiLKYN0b7MHSyef2akVwMUiozokObc6BgYrMsCxuDWdRrxcWe8U02rnmaCMTNFd6xg5+mh6Hd/t1Zyc/PUT26fmxvP8Y
80s1u2OqHYTm0Fd/2Mp/6JgP9Z1TR9ASm2PyzxXsHLQKjsoaCsSWhgreJsjDWjWSba/V9refaFQlYDw/k4kYt92tpXxQbPiMK+5l7Hf9Oea2He3yq1g2u9JA5g+x5L+y
DiC5mkoPFHEU8Y/jMM9bLXmXi0cBBNzIp1U7i75hqCAPwu3/KS3b5q1rsUYSHUBt/dkT9ixZTJf4w6+0TRNpg+eyjcHGEigc7zLy/sRJUIlv90RRDf67G3YUVjVlvZ3B
LP+fkGk1qObC/MHRAAOxW+JGL+fhYbZ6K1gZzzIHUh3cD8dBQBgcZjBz164qcx/8savNdR6LNsDp6j4l297kbVZqk5Dk5jsxZ+awdOF5hxJIVSkI7KbAY9btSsWgi6RQ
cDPp/9zjOlRzwTLFveh9SvGrnng6Zun0R29Zp9mK2L/sAasrrYd9Fjb4aXGdu1pdRU7c4+AcsoCp8kKEqxqyMqaQEYVFssLMtkjFCl4yvaXKiCbRJr2HgYyrX3ljAm2I
ncBbaCvUZbZ0R3BeM75ZSltdDv0yE3byUoH/sNuz/KcN4FjMenpr0KQRNWEPS1m7yogm0Sa9h4GMq195YwJtiBJGqJWn1t/qGroimMFAGFYr3JLpGcmtgQ2/Aek+GcDL
yogm0Sa9h4GMq195YwJtiLziLrYXES/CFG1ZCH1SN2XUoJ8AZNRb3Haez7R21PWvl0mjURa8u6sIGUa7IOUHDcqIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKod
PfM57ZQJ1+rjDf/0jWoaisqIJtEmvYeBjKtfeWMCbYisD+Mswa+YZU19VKqRMUbvH+SKzx728+3vqrjqrX+uNkAUo6urhPISUsowl/2BdGzKiCbRJr2HgYyrX3ljAm2I
FdJkT329i7COnhM1KYxKoTYHXYgL+ycDuhVAjc2Hz249byeZFLWBz5MiOduS6koFvV8gaMhEQEQ6/OIyj+neUrVjndZ97K9Ai+1BkPzcyuiVjwyx4rk7hBA3iByP1ZoC
cmNCpBnjWbsQW9+auUYlAapdTQe1P54xVOX2gkGNl9fgedcEGRbG60c1ea5TcACkYAyEzu4aubwXNbGVPKkCDCrwJ30n5KU677EG5Q/JndwEdB4SCYWlTZXahmtbyiu0
V1oe5Eu5r/e1l98li149BcLyT3RKeBcg+5fDaYawF8RAyaqwkAgzq4ApJkwTRqQMsqX9wTkWfLIFmYB2lI8EoUR5fAOqRMZI8caN1bbRFZXb9mVCyX6YOPucAu5kGysn
+D0HgtFKzfcPpnHgjrHhMO0uEXmWTy1Uj4Sehymt/kka//rs0DUYqzgIWeK09g5oia9fmNFgGjI/5LT99C91Gp6tFhKLAQFqkrN6RqgFI5vdnFF/pAXdg6FdAIyt1HS9
3dghmcK1x9mAo5MAj5zqzIICtUaXATIf11KzYbAa453DDkBpMMMuC3aEyxQL/uJA071Ryi+qiA0Hhdug1eNnNn1IKEo2SdJnyzr0362qFc5X28+4p49lSLsvpCISJXvN
i2Brb2P1bNYdqcrS0QfexBSNyUk5VeZ7+SqbWWfc3KKJ4+W0Fr4xEjv8T/zSik94coAjxvjxhUb5Otvh+49Oz8qIJtEmvYeBjKtfeWMCbYjpx1X7c42EOenspv0DO9xC
6AlCf8lzwqQQqd16Lrsd33DvRSfVD0hRzob3Uax5dcCSyv7mlCuiNFcSWG5SSuJgVovpwjX66oeTMs7V+XIbqC9xql7ws+8iYnKT35aZ2tAy4cZoWKoLRVrjQc52GLJL
nkPELMSQBI3KYVRngPExRkKxBbmrgyEq1mtJcdiOLOfXJ4ps8BDtBhJsiekfumSSQsdjCaTmfg/wrR+cdLwJGW3DGzAHATFJyRAQ8K0kHAJcxEYlu0KnEwuTZqDMyJSG
yogm0Sa9h4GMq195YwJtiDZlloNdhddpYOAaTVdVPMcr+2eaYlBnTWBxbOnmNWO9yZE8d/Myari4nkWYlJSDYb0lSLUI6L+4GCIkVAznFYMH+NW1NjHrI5s9sTqw6elF
T3uOYf81ndVatzKlsfwFeT1vJ5kUtYHPkyI525LqSgWDcRdOfnzDCIY08vsxLu17jdJCa+YLMQbsRqV/7VaoHf5Y0IrBpttDMmPH6IkfPmgjn1Uzj5jYW4gP/IcOKkoR
27JEuq2bwMWufo6wQU97nAFWJ4YrzczUJzWRf+tmTYNgDITO7hq5vBc1sZU8qQIMcgcuqXz8VKFxDjVJUfNjdgYBZKGW20y0NuyBLre4D5GKq59VLpM5SEI2mM4luCdO
GcEA1RzHrVjxmyxb/aN5Zh+A6OV2z+UESB0Wf+AS/jnO+WSuEazdF2wIzgboayUUkoMB2n9gv14Fx8cHb04jDjTecjcMHpjW28W8vTOGKM+SNw09cGng8UC0zuarcnzV
7RJb/9kOnvUS7RTAWpVh1IU5cdRuF9j/DbP54eKnvCfP6WTxGYatyFwk/zfK4u5zS2DiPrjaI13r0PaE+NA958U02rnmaCMTNFd6xg5+mh7J+XumzoWseXbWErxMkB/y
PBMoSA+R/4beemn/L1nqhTk5eTLEg2GNphNUI+ilb2+UVNyq2AQPD9kvJB4JjOspUMdul97V65UXqWOwmzgR4uj6Lraqu9zXKuFhmlQpl1O2He3yq1g2u9JA5g+x5L+y
CQQ7ZF/uGF3uJggWJ63kECtPQgGgvhnT6E6HCAMb+XjvE2x9KdrA+nTjXyN2og9Ycjrg2djo1TimXlYnaDFobHY3cu4OEnYJiwLELIV8Fw6iz/T6Tk7W4zOuo34YRfeK
LP+fkGk1qObC/MHRAAOxW0XcuT70YJa8HUi/mkxwtk1uE8JomAdCaF3g9Zf84UgZSB6jnxB7C06R0m4uR2cisgIP5RvZNy6IzJlWXrB9736dwFtoK9RltnRHcF4zvllK
aVpDSJEedvgdZYNODD1MofGrnng6Zun0R29Zp9mK2L/sAasrrYd9Fjb4aXGdu1pdEkaolafW3+oauiKYwUAYVtlvEaIkTB8kzut4GGcFD7TKiCbRJr2HgYyrX3ljAm2I
36XbMRKQePRpdT6uwSSooRT5woCDkTCoNf17S+G9NfEIIiFhh/rwGi/cIwrDjvohyogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh3aq9oCstI3szuEOn3CsVOA
yogm0Sa9h4GMq195YwJtiKwP4yzBr5hlTX1UqpExRu939ESXTnGGSzLJD2Jvh67Fl0mjURa8u6sIGUa7IOUHDcqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqh
EFft8SMztCcFDEPYx5CHHsqIJtEmvYeBjKtfeWMCbYi9XyBoyERARDr84jKP6d5SH3ztotOdSpTlYENLFvACxya+ATwoO4W/MoO0lSRGkf3KiCbRJr2HgYyrX3ljAm2I
0vZ/C5D4uxV8hGR06yAxc+pKep3K4KKr1fcrHssd1vxcNTOtCc+GcEoyWXd2sbjuKvAnfSfkpTrvsQblD8md3MHGuSRZBeQ1QlxYdvj3E5jcTVU8qyXCSTScAfytCAo1
M+rZT0ajHz7sixcQqGUHA/a7MB+UZd1JHic/n+t60+8GpBi/ZlTQ+Ls+seMWoFIFp96W3VtnIC3fvWoipO87Qtv2ZULJfpg4+5wC7mQbKycsxfQP0ynhZvZkYjfJGIne
nxxh1l6Uk6O89GaCSLA9NDelwudn1uXM+2+tqQjKdgMpsBaa+693yKVXWJwNX13L2kFFbNZri1cSG4AU5NQQjmmE12LHyNDpAezjzvuWTsjd2CGZwrXH2YCjkwCPnOrM
RVZgZ4SUeZDIi/ol/+xkwY3WUseYTOJjnm586pqEQkyCAe9FCVw54ZhuZT1+mcPjgRrInBgZD19HN9j5BZzno0h22QhKHYp9svQ1K+BB1hcGjK2ckCWSEBRoke9aL+NG
FI3JSTlV5nv5KptZZ9zcooBdu1pYhLd6VJjo2l0Ps9sPOamloz5qDX0bZ2StwcDfoaXMr+7DukL/82T9ck0fwDg+w3aQGvSEU5mfr0QFNNDXWqgUmTx4guBJbDM7pxvs
ouQU9H5luGUgxrLFEfdAxqP4K3Cg89Rtl0fmHCVx4N5NW8suQB1EvYjwuk7vCF78QPi+gV8w7hvjt+xCPl/2XV9J9A7WityQch1s0PeddJxyBy6pfPxUoXEONUlR82N2
hyEg5O8ocddmcD5vnDnXu4G11pEGp45MPlRTPL7gr4BkY9y34BxWEvtb/WwWkMBafZ2IxyvvRO+2K4Lu9BD75t4ER6ENG7m0FDD1bgBFTDqsuvWuSn8ecEZ0VfEJOOCq
hQwNEm/Coz7kgqDyAPzL0qwjK3BzueTz55ezm5Vm7pMDqOkDIyv7RHxfx/5zrs567CIc84HygzArxiUWOLGZGAcmGxct8u9B2WKVHZWZinWQxqeAvLOlVwcrs619CcDe
SZXdRwN4saED/s81w/rdTAcIGKSnElmvLInZ9BdAcmHKiCbRJr2HgYyrX3ljAm2I9rswH5Rl3UkeJz+f63rT72wIx7W1IxuzCcIi33W0JFyLYGtvY/Vs1h2pytLRB97E
vTr8Pu0EBlSSjvHbxZ0KKCHVmJK/R5yzU4vUoGAcMyegU3uAd5P5mx4yFH6qOu0i6oYqzNSVUKvxKjQcQIK+87j0ZFLMbeTSEiSVpuidBlBFl9LipQMwTP0E/gMuXhd1
pWrYDxMY8EpFGcqFD12gzra3ETb7Tqgze5LTRAo79P1h8mDhJ46N/Y2DEtDyryGTvtU0Bj4uTOQNJyq1bemFyLynG8KyleKT9T08jl1zlLUJ+zj9Zc/hZq8MCTh0LiPr
T0AdSo0+Ioxd3pOapgecMQyV8DmAK9BvtGj9B2MSMcMTvLvRRbSkEV2Cn+ID+F/4ZBW6B8WbMtfByuI0e1tCQNOv0ql5LTwWyRSKRdMk84nKiCbRJr2HgYyrX3ljAm2I
Msq5IlJVpr6vp3TahhcLfsM6KtTMBc1app+Bscgh1EDJCofg9yt2CUjfM6ZEu6U+ClCZ7L848VXrkTThzV+hlYP4KgKvHDh+lxGjf3WV1jjS9n8LkPi7FXyEZHTrIDFz
YU4xmip9A9N+SeERW2GIDLJ7D5gopf3ltziTucnB4wqmCTMrxQsCGtgx/j+OC1/V01JX1VJmBM3Mqo7dye/6hi3EKpEm2wIjPE/+XdSodx52A5eCU4/6N2w/Xr2Pmeo1
LmKRiI2lIu7X97POMWrj6xTpJIAL0xPlDIsMt5oW9ZeGqYElDOrGcWykCVdW2hGHSVnapmS7/B24/ISf4QIBq/5q//qpyStb3Rvrd5jFSMyLYGtvY/Vs1h2pytLRB97E
SdQXT+AQ2BgoYmC91QBgpEb7a4HmOPojlRitOEVQ45DTIZGc9kTWzrYMDyDvnYgc/GzqDjB5zK2c6GwB5P9jobj0ZFLMbeTSEiSVpuidBlC4tSXd6xGN3Z65u8uMhtDq
lwXySC2tKy32yeglXMcWP8qIJtEmvYeBjKtfeWMCbYgsGYz5CqUEgo522DU+NNCcw227VC4DMoLGHecuttu6U1rk1RUIu2pRBpMw81Ln+L6eqts76WOv9BASMXPcGYV3
UBThsQjmS0ur+XHUzMZ5k6VXd83dOClpLQ+xdIQvkcbrdjvpQvbHmsSDDXbKQ7pfyogm0Sa9h4GMq195YwJtiAfMz+29hT6raoFciUGFaZRa9JeJrlpd4HBOrfnQXdNi
ia9fmNFgGjI/5LT99C91GmeNmc8gsyIKYoOinUJT8pTKiCbRJr2HgYyrX3ljAm2ITHP/CyloxbBdUvKssKHJddp8KaxIxCfwRJJPZaJ4EimeQ8QsxJAEjcphVGeA8TFG
/mkRXqoMjGUEX+4YTuPUZLJ7D5gopf3ltziTucnB4wr19eswn9HLHt1MO1f6Mv3vA/1sSabum0a5+IQ7CMWTSogkScrPGn2suDPtYWT77jpvyk7qfn/TI+80VrKqPGG7
LpIc/SRxK5iEqxNSsQy0fKWK9z3JeXEpLP2cG6iw28a/PAw8cqiFYEmrXInGx+Le3gRHoQ0bubQUMPVuAEVMOidbYelD9SeuhtTOn320HTfWfvqzV2nuF8JLgwlFrZ10
rCMrcHO55PPnl7OblWbuk5SyMCv1xV8A4+uF2Ip+nRLd93Jg0pPUijZXofrfCAqhqU6BLDyPrES+eY49ZMLZemnOaypUlqFhFnm5npN8gtNJld1HA3ixoQP+zzXD+t1M
QBFHEpMkmNjE0KTyVEAsWDLhxmhYqgtFWuNBznYYskv2uzAflGXdSR4nP5/retPvgyLX9sw8mdwB9/kJkX5jN8qIJtEmvYeBjKtfeWMCbYj0FcrNa6/DHKdR42sEUCkf
dbhNMq13WxIV1kkcCXys8enHVftzjYQ56eym/QM73EI4hDZrmAdYQWC+Rdt4rrb2QeB647ENxuW+M2jSpBNlUkWX0uKlAzBM/QT+Ay5eF3UX04s7GpOWe+lBsEcIH590
9PuGTLwaVy16jpBhbuww1D0JrlFHTB1AKW1s/+7AKB0KjsoaCsSWhgreJsjDWjWS84TlkgEpyli/8oSmxFQMQW8niTk+7ruB/WWlZ23Zah6CnmmjWbEdLVCw0xnGsVND
6BOBKiCxk5N620kFEkkFxdY+gf/RVaKibyXFhff5cgrgRttzmwLZ+nQjtyw1AL2Vheos7k708fsiWcjmgeuLJcULTu87YwhicITWZpK0O9JMa+7PbL4Frz6E7z4XCFQ6
Q79gZVwpLWS+ToQlDhqj/GscVRQbuNSp17eIXJI5C0+tG5/mT54mfrRn6WGa2XwxXDaoZUqFYDT9k7bC46uTL6pdTQe1P54xVOX2gkGNl9dPD8oXvcFTL1IBfux5TpYB
yogm0Sa9h4GMq195YwJtiFKCG2Baz0Az0gGbyqCdyyokF9dvoI2mAgTUeUHLCVdIfUgoSjZJ0mfLOvTfraoVzpWAhC8cTeyxMA5fKRcM2CdNf3RUCPmzaE3QNwrVymL0
krjwBupVPJps1DrYrrTvQMqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iqcUqjgFWNX7Q3iT+5ZG8XT5RU3KrYBA8P2S8kHgmM6yljyA49B8xLBgvQIkybRuzT
10+KIXsFYTOG6b0aut2at8YrrLBxLv2TQGxj8BkGeNJUvdyI2iZhAYK9QgCipoLxhqfJbKCQXHya2CB70Q7cI8W0UEnsETxRX4aK5P5x6x6Iw7HTqRSK+lmh0QgwU4FN
yogm0Sa9h4GMq195YwJtiMOg4wWodBrNnglhNjQgX/4GgyIc/DkbJJinnUgBuzjB+xhd4ZFcymQKDOaSRoNR70wAmsMeYpW4YWfGoZsD/WnKiCbRJr2HgYyrX3ljAm2I
nRaX03aQ7Emu1LPCy5ShPCEjbEjQ8i1SC8ooJ4dR9jPKiCbRJr2HgYyrX3ljAm2Il4o3ttizpWWaoxKVK+bDJMqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
SrPcvLPYyFjjYiFT9IiUB0GXpZXyFfkhDGEWD774oi9ErsYoRPN1Cw1jbTE+NyhEXNMhCHymiiPp+OD9jGHFtbIT4SXjgq8NNwI9BCre4Q61LHd36Oay4i7slx7SJoaR
sT8Bs0NZZ8sGO61iBtfwG3FsgSwKI7PGeEPmnWTgkf+Li8tZT59+8lnmoiK10Vdii2Brb2P1bNYdqcrS0QfexGPIDj0HzEsGC9AiTJtG7NPIhhD76vmdN72p1ECVhN29
yogm0Sa9h4GMq195YwJtiNMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/opZGcqEr4VEXxRwAihCVK8Frk1RUIu2pRBpMw81Ln+L4fx5Jb2INXjs1+ZGD2snZ4
iMwH3NDvlqUs/QTvk0wTLcqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqhgHU6tMXhWGtdTKOKVdJ4IMqIJtEmvYeBjKtfeWMCbYgbnAXdZ4PD7Q6ReHlONAYL
1yeKbPAQ7QYSbInpH7pkksqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFGAkzUKh+ZI77hc6HeH6sjhYCmNxzirTYd7fXcs4sXVIRSeTJhE45qmN8ZpsAfXCcV
4xFg9IsPGABCFjL60MwXA19+MMqNYVnbPVQwWtV+vgreBEehDRu5tBQw9W4ARUw63A/HQUAYHGYwc9euKnMf/Ky7AieKG2XhjDpp8/u2lNePRT4yVnQygGoejnW031O6
btTcjOX8MrrDhgB5lsMKvJCD7qAhAHIHQ2KxQHxrQacyzpinzexsSKNI9UWW2xEw9rswH5Rl3UkeJz+f63rT77111QhUeY0Vt/OTOatyTvPAOKM8gFdujXkrsIGWPG9g
XZpyYW+WQ+Y4dri3SmpzUJ/5JZYlSzIWeUYgMrSqKrT8mRtJCSknap5v+hx+YwJRg3EXTn58wwiGNPL7MS7te1SC4Ivaba+mMnZsrN6XPMCXGEFER09NLos2DtV4QrWk
4Ebbc5sC2fp0I7csNQC9leSRjv0GsO4AXU3qKeON0XkBOlMYr4/5DVlh1mkSMGibyogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YXLum6X9JKMqRIWmkykCsmc
rl6GzEjFrToJhl3WfxMF9265XqCu308jQ3yWo6+pBTsiXU29vnudd/I3rR27Uijobj3Ko4+CjH8yg9uuGxmZnYEayJwYGQ9fRzfY+QWc56OjaqOmB8Gbu+bzvDlR+Fdz
BoytnJAlkhAUaJHvWi/jRmPIDj0HzEsGC9AiTJtG7NPzj+K8TMdkjDnDU9uCZ1CVUEsa4O3+p+CZ++chvFma0NMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o
DeBYzHp6a9CkETVhD0tZu1rk1RUIu2pRBpMw81Ln+L4fx5Jb2INXjs1+ZGD2snZ4nSMu4njndQX2wMg4Enhkk8qIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqh
K/Y4Zumu/OIywkYyUMV5n8qIJtEmvYeBjKtfeWMCbYg2vA7A1pFw33FVfP3pDs+0XIA6IN7aK96lFqPI7XaeZsqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFG
26IIS3M7uttdAWjIqnti5dcnimzwEO0GEmyJ6R+6ZJJSeTJhE45qmN8ZpsAfXCcVz/SQRObbKQHuPZovcLPE+r7GHktMUlHHsWDlTchce0jeBEehDRu5tBQw9W4ARUw6
K09CAaC+GdPoTocIAxv5eLYEu5VV6RvRfKX0i2y39rtgRjsBpYUIdhlxC9oFNuSNW+XiRD9/2CvFZMe9oOrJY43WUseYTOJjnm586pqEQkw0lxWeXycLaUmdrNjuO0/Z
QMmqsJAIM6uAKSZME0akDB6IukAjWr7fhkSotD+/bpCkx2S+Dhp49npnR7LPDRwiyDZ/MjIBmTwQZtMW8xLfa8KlVFlFIY4fc3p6N/DrPFK2He3yq1g2u9JA5g+x5L+y
PSN7k7iGlVp8dbcQNm9I8nwuCEegFy4Sxost61XiCXRlL14oNYYl8oQ4/eLCFWb4jHuTCHrDuYMD1aHwijEX1F+7Kdz0gey5ty980iI1A/u2BLuVVekb0Xyl9Itst/a7
bZq+2OTrgHGsUp66ydkjExJGqJWn1t/qGroimMFAGFbie1gOmy8QAJbGvaXIBYsRyogm0Sa9h4GMq195YwJtiB0mmPTpDtYNHPj7jwGt5kOEuTXwTF+5N0QgHEzjq7Z7
i2Brb2P1bNYdqcrS0QfexH1IKEo2SdJnyzr0362qFc7z9LzmHRLYi24tLMnDcOeDXIA6IN7aK96lFqPI7XaeZpTwVTaMGH0aC+klaOr3Y2jDOjZkUNt07xV/OvkF6rgM
zokdfAWKlXjJHMWLsHayodMhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbgugSHUx0t1kAEhXJrUNlTrVrk1RUIu2pRBpMw81Ln+L4fx5Jb2INXjs1+ZGD2snZ4
EILQMUa8rQzw27FOlL6t8MqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqhxV32myuZPEAw4C+6VVBiT6felt1bZyAt371qIqTvO0Ki/jXXpo7RDQkl3aP2X67b
cGR4YExAy2v3hbu5mfwmxICmNxzirTYd7fXcs4sXVIShjhkW0xZR4jr1EKYyTILNQdnUzwo50ypcHRGtXiihEWTjwZHrTCzECRZLp2toLUHCcIXytZGh9mZs4aJ9+ttM
ZBbR0W07Xq/msFxe7OI4KpgP9Z1TR9ASm2PyzxXsHLQTnnY3PaLBCp8wR3PX8eJ0K09CAaC+GdPoTocIAxv5eEohNJtNgnDVEe/C9LawVURySeWx2QsTJ8dDZ4L5/5PZ
W+XiRD9/2CvFZMe9oOrJY4mn0fTXKRFN5DZgpLIwN8bdBK86ougUBevUt2vBNSPKpSbIbr2pScoRwKyIYeaPVHyM2VdxhFbJxFDohtd3+ehEeXwDqkTGSPHGjdW20RWV
yDZ/MjIBmTwQZtMW8xLfa4fi37CEzPd2G6nTl+T4wxqXGEFER09NLos2DtV4QrWk9PuGTLwaVy16jpBhbuww1CQ6rCycCPutlY134NJEJVNfKzomxJ1htltGnRRtNUv4
3GVHMZKHzskyz5psPuSBy1+7Kdz0gey5ty980iI1A/tKITSbTYJw1RHvwvS2sFVEI8XZSVq+8r3SwyDHpQhuOhJGqJWn1t/qGroimMFAGFZp1g6IvjjF5ujEXdOtLd1x
071Ryi+qiA0Hhdug1eNnNh0mmPTpDtYNHPj7jwGt5kPwt8wXbtO8H7oglc9ISu0FBoytnJAlkhAUaJHvWi/jRn1IKEo2SdJnyzr0362qFc7fmJUvxTrfa3xhLFsYZoFi
2nwprEjEJ/BEkk9longSKZTwVTaMGH0aC+klaOr3Y2jDOjZkUNt07xV/OvkF6rgMSJhpOFU3JEBDrxHqs9QEr9MhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbg
jnu3S4H1Oil4ozRsf7pk71rk1RUIu2pRBpMw81Ln+L4fx5Jb2INXjs1+ZGD2snZ4u6KnBTD1tZKd1IQeR3i0wsqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqh
4wlF7+cGjzD7nnZFThs7Ay5ikYiNpSLu1/ezzjFq4+tLVUG8+Ktjg9zMamTHAuxnBONagr2PcZ9zXBKBZWw6OVSdgNgb30eMafXQXIQNIFyeQ8QsxJAEjcphVGeA8TFG
wb2D1vR89jzRB3iMn2RtHeSlV3P8KTsnpYOsGxat/XaRptehNO/fVB4PS8KB2zenHNfuQvYsDCb1r0BdkJ0NGsc40kxf+lZn34bO1gpWUTv3H0C0h8QulsHEaT5tT232
3A/HQUAYHGYwc9euKnMf/P7yMDK937qwFptBMWi4eR/1/+JSoPeO87xFaG6zYYtqAMdxpH2heDRRpKcBwQbDYYAUdFsHC3k6TqDkWxf/3mYEWzcW8X/s/esqwkM0mpq/
9rswH5Rl3UkeJz+f63rT7427HLN6Tqs86gIB+9BtPAoGjK2ckCWSEBRoke9aL+NGcR5GzyiEvYh/W4npYbxrXzKekqoS9XbNXaa4PnNodBmpke42a8avDa8r8kKYOYu9
HxD25uf2vH7yOSe3Uar9PZMEygrQ9+FtWyjlwNGLxA8lC26/jOtjVne7S7jcGXJphrvlEegmBpYWByI/lIPadw54gSc973VzN8T40a4nxGI8rQ/H+Chw6MmitXJ91FsC
7P7kec8cXWBcdxverVThJiqPZvSsJfn1fRBz/Evb+4olusyZNLKP2f5DvCNO16FacoAjxvjxhUb5Otvh+49Oz8qIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17
VILgi9ptr6Yydmys3pc8wH1mwD3CEYtXA4GZ7WwI/NDkInEXnwPC4/4rNc3ldMDDyHfX90Etu+C/RxWSmaPQ8shh1ljxbJsNGeMW9WN4kZFcgDog3tor3qUWo8jtdp5m
6cdV+3ONhDnp7Kb9AzvcQnrL2LfQr3s4seH0/fcu7yVUnYDYG99HjGn10FyEDSBc0P1z7btnOqj0MScDpSTFynHgZxQnts2mIRKhpHF9sqUGRBvgNgk4nZQd8LxzLf2y
yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60++9ddUIVHmNFbfzkzmrck7zp96W3VtnIC3fvWoipO87QgFuetFy/TYk9EoJGmyb8NCMd+0Q4S2bwbxGzPLLl0dG
gKY3HOKtNh3t9dyzixdUhMqIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKodDGGjYSX/mJhUZdMFPwZj1svEocG2y9PWWO1ABPG9Fko1O9BFyh+oKBE8Rum4OZBp
3f8zqqknTv3zUOe2z0/xCJDF+xfu4ZNyscJBSqfM92AJBDtkX+4YXe4mCBYnreQQ3A/HQUAYHGYwc9euKnMf/Ky7AieKG2XhjDpp8/u2lNemxQcg1wpsOVNIwDoOCCoL
SarFW1S7xkQMidlrgHnCjxV2EeptmemmdGcA/qS/vtz31qy+VPwjRFqTJ6z2aHYxcgcuqXz8VKFxDjVJUfNjdkT0lZagVCqYs/29yaA+ICAjoxk4n4lTuIuj7F1RIGUS
xDi6C0SS8eYFRnmQEJGlhiIEBeGptREpFM4lDaupomlIHqOfEHsLTpHSbi5HZyKy3W0mzfqhJn+IHnJip+g2dJ5DxCzEkASNymFUZ4DxMUYCTNQqH5kjvuFzod4fqyOF
sECBbdgdd4Jyfk9VZ2LW+OKStgkrZ629oZbxnB8ICv8lbhvTqd1bl/DXCTVU2mzWXys6JsSdYbZbRp0UbTVL+EtEfLMsbBfii5nOjdUXRfMpsBaa+693yKVXWJwNX13L
satE87EvVlmGcqF1u9dvhsZYsRGgBt5FiwE6FcJmjRvHZphWbz6AyKF1K1Ld2iG/YYgRE/wAiEQRpVw3FFd3SGC97zKY2QP3jtmg5o7+vAUWiP6smxOZ1pZWxVkIHXV7
dEMpVk0/iVLB/Xc8gKO+A+T/ohkl0SN5+FwdXSNiFiDKiCbRJr2HgYyrX3ljAm2IooQOPG3OcfrPF0EFXlE0dgi9JRYLPs8uhpFWo8kbyAKdIy7ieOd1BfbAyDgSeGST
yogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBlJBcl1lTcVejt778Q1XBJIyogm0Sa9h4GMq195YwJtiOGGDY495tU//ZFkpKIypcvwvDHFyk3aI4WgeFu1/yEq
2IxgPx4X0/eBdEw8eySRiNMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/ovsYeS0xSUcexYOVNyFx7SPDuFpFTYUg8RVN19ERnN4udX5W7Jzi7Wh08kCgAzZzq
Rpj/0IKCZOn8728fCke7+05Cr2ncmGPf3ZyQ3B3aJYk2ZZaDXYXXaWDgGk1XVTzHlrG/uQOgf8kAh5goiNIaoGoFHXu1ZCmG3bhV3wbEcCEXOKIoyZHj/kcU+FeB2LVw
BStOHwZg8x9iM7M4icetBRBngsnIfRnQs0QWNrmeMHRxU0NIHL16r5NXe09sJLq3fUgoSjZJ0mfLOvTfraoVzhoZ5pG2DAwVL0uITmd2OLZEeXwDqkTGSPHGjdW20RWV
hMhbM9s0YrP3aHIgmqJs/QLqHGXEYhCfbIHG7y1d2rarcuzjLW7FpvhiGZ/1j4fdLCt+lDet2RSaOErQw1fZy3iCUkzMYCZ+Pgy0vo+tE1NHLkFi/FVFijqlfbdHCCXX
oaXMr+7DukL/82T9ck0fwFQ+EJ4gyq0D07Q0/RTPhWhd383aHFG8pLoRz/CmKgF1nxxh1l6Uk6O89GaCSLA9NFtC1sTHSlKTj4dIga3WzeMSRqiVp9bf6hq6IpjBQBhW
Vp2lCnu6UobJcc5iztrUg8qIJtEmvYeBjKtfeWMCbYhJtbgU+uAcoZXR8mGuIlTVbTGiGNLNGzy2EsRf7D6gf18ii/3q5rc5+VzljPNgB0NPQB1KjT4ijF3ek5qmB5wx
PBMoSA+R/4beemn/L1nqhbxmOdu4zwByVpPCS0UvMp0qj2b0rCX59X0Qc/xL2/uKPTCOW0L6tA0RU/Uqf982LkASBELQXIlPfpRcs5I9LSyojOXOHf9/aPv8yX+Q/DW2
g3EXTn58wwiGNPL7MS7te/aWoKegf41mbGTwL6/1N9lZV6FrtVlhP2ePcYaM6oyU5CJxF58DwuP+KzXN5XTAw8h31/dBLbvgv0cVkpmj0PJI1mh1FNCh8htDhUnJ/pgZ
EeC7kPmsKMQZKsAumoli9+nHVftzjYQ56eym/QM73EKiLtgP+Sx0MbomDLBjh0VFrz6jMcSqW3uL12h3c5iq49sSlW1oJVb7P0LpuQJagLY6RWlfWY8ltLyghV5d4B9v
rE8w/B0dn3x9B3SGQiZdjGaVJIJtmjFj+Xv6fpVoy0RAyaqwkAgzq4ApJkwTRqQMS9nYgO0pBt2d99Nl/fK+st7YN+iWSI0zfA+1UPUf1bLL4o8/2IkGAXivjsMiLlEG
HtJLa4LCBk/QpJrL5CdRIVAQ1lbBQAuFS5P0/H1BpgbYlKH5QpEow+woh2/lKSwmHnxxE58x7qzsr23/eeD5yt8/mFB+bRSgqpsPMQv7+KvKiCbRJr2HgYyrX3ljAm2I
lWY9F+C/hIS5f8jz1U2I4jSxPFJzcVv4lAwB0CeOj8nl86uJw5gW1jrjD4MYUNRdksVCEwYQqdTtxoDIQbz5HStPQgGgvhnT6E6HCAMb+Xgl1Awz63XoW5yxuRAhSpt0
SZXdRwN4saED/s81w/rdTAqJrloSNP0zFCLM92m3MQCHz51KHGIS3SUHm6DHEstpNbCE3UIUUabPsEYLmtQL03IHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+R
drPSVDp4R4N+iUp6b203Po7iQ7nBaKh+iDx0aaXgHgAxsUfkMkvKO8mmX6YN8HXiBobYEQ+Nh06EWNOfSwHiY9g983Hn8j/ZAnJmjZA+dHmhjhkW0xZR4jr1EKYyTILN
coEKfG6UnScpy/Zq0Z3c+Ytga29j9WzWHanK0tEH3sRA24bVgXQMxBqg+LqBsqdysNzzuRNBnsXJuVOgboO8mpcKBHhjfFtwMzdJuGYXGe/7rICpy6vrQuFpgCGDT3b1
ia9fmNFgGjI/5LT99C91GmDL2lFb4D3O0vJoHJ8YD+nYjGA/HhfT94F0TDx7JJGI0iOvNx8yGsuBUNl6SE4EbH1FKE5fikB3n8aah826wa/0Tfi2EqWlM8kxQQH67xAE
yogm0Sa9h4GMq195YwJtiHRDKVZNP4lSwf13PICjvgOH8A+0ic+UARkcf+OWHljXyogm0Sa9h4GMq195YwJtiKKEDjxtznH6zxdBBV5RNHYIvSUWCz7PLoaRVqPJG8gC
UYmdmNljiQ0Nt83avCJ0DFTGlDJ3QcBfpMDJLF74XkZuE8JomAdCaF3g9Zf84UgZPIv3esxXs81bY9Heho67AMqIJtEmvYeBjKtfeWMCbYgfW3in/VVDt0p2sjJRBn50
IAfFXjDjb8IaS693+SRdxiM911KnflKdPBdpxJANGWnTIZGc9kTWzrYMDyDvnYgckjcNPXBp4PFAtM7mq3J81RjeYSm2VM34dabATX+7JjHw7haRU2FIPEVTdfREZzeL
nV+Vuyc4u1odPJAoAM2c6llY5rgea9KyOtkQSzEckV7XJ4ps8BDtBhJsiekfumSSNmWWg12F12lg4BpNV1U8x5G4hFclJcRLbxcCqfx48y/d93Jg0pPUijZXofrfCAqh
bZoZm0kBbv+EGdyEIDGEOLac7MX0YFQB9C70AlP0sdeDzO2laKku+IzbkLNqgNt1+6yAqcur60LhaYAhg0929YEayJwYGQ9fRzfY+QWc56N1Xr5Sm4WWlwl/Bh4RU9Wy
MuHGaFiqC0Va40HOdhiyS4TIWzPbNGKz92hyIJqibP0C6hxlxGIQn2yBxu8tXdq21aN4TXcq8iYXu7plxrx41cqIJtEmvYeBjKtfeWMCbYiqXU0HtT+eMVTl9oJBjZfX
q+Ojthg7dKHBO3DcOzPliBYxVqT8lByLUn8UlLTREaM92E4S/6aE1yRdKhgBsVYi/cORsL++nfNhMApynjsK41WVXdPRucqNdCNmtv0wgS3j8Ei39Tc1oKpr3Yw9evoZ
bcx9A3euJafUPZh7l1vZhTkUon54Mw0hiSb15VyZJN7KiCbRJr2HgYyrX3ljAm2IgnVXWJdrlpoWPt54kYLtFg5pQuUrhjkblzQeOns6JP5rBWhxdvrZJ8ZSPEokRQUA
T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCBtjiFJkmFARR3dxerGQWiLKo9m9Kwl+fV9EHP8S9v7iuSK3BoZ1PvdzYR5cTCKabILMDWCIBP1+IpSQi+0s7Gq
nZmsuqL6lQq2Rh+X/W+b9YNxF05+fMMIhjTy+zEu7XvaxJ5t5YtgAOVeB5hK7WrB8FpnaOU8oOxbgtDgG8ilO+QicRefA8Lj/is1zeV0wMORpQjoF0MHhwFqQCq8NNbS
idfNdOBNVaHjqjsPhxif5C536WTFDIpNI7Bv8oKTuB2gU3uAd5P5mx4yFH6qOu0ixv2gh85QdGJLxa2MGvWJGNjGYyvp/mIbJmfNVRQ8DTDbEpVtaCVW+z9C6bkCWoC2
1kDeTQSet2EUifMY1sn83AhvAbk1s4BnjpVBYGW1nPBjiyjfzVTPXrFbZ99I+uLJ9rswH5Rl3UkeJz+f63rT76zmEvI8lYdwX86vIAnP9JHKiCbRJr2HgYyrX3ljAm2I
dtP9lUIO57/l3EXRUcfl/GdyQjWL9s7MOjuGNxYddacPZL2lz+T0HMwj+3hkCNgZyogm0Sa9h4GMq195YwJtiIRzeYR/RfNl5UciUvKeH6VMAJrDHmKVuGFnxqGbA/1p
yogm0Sa9h4GMq195YwJtiC7UEwkjnGxYq+DD7vjTLkbKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiN4ER6ENG7m0FDD1bgBFTDrNXtLtfDARzwmVP2fLjDqL
yfD4Ai82Av1anYKXUvVrL0mV3UcDeLGhA/7PNcP63UwuyHpldRj3E3yXLr4oDIO+yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhCIf7qwLt9U+/9lG2X0qvj
q5S1ajz0CkT5Q/7n0vfFD57OCiMGcKZ+kbnsuetQ//KQGRB/j25c0O1QYk/jJYA6lEZaxz3AupFYYRz6UalYyRBV1Hzn7iNe66/pbDVS+Q3NK1L3pvXcN6PGuMClU621
qK6l3ShblWWNIdaLHPMuUqmxGTVOugBbfQ/emIGXZhxyBy6pfPxUoXEONUlR82N2jzyH6XoYf6CqDONvEXdhfKP0a7wATdnuiWFRXeN9NBSEyFsz2zRis/dociCaomz9
QeIhi6jhngAy42zoY4nkuFjDFh5JMDb2TZSH5Rx8vJF9SChKNknSZ8s69N+tqhXOvKKaQDraTz2M1IAHG7UZA7yWYnGvLSbIxq+ET/7rIK+Mb/a7iO5xuloQcxWXFwIN
4OVTuhYBZ1AC/Pdv+X5t62OLKN/NVM9esVtn30j64snnUrwFTsoIgYnw11fU3eejiwc5SVXENxHa/L7mqET3LHN+WqvorE84iDJuOp9s+0WDZTYf+QvAwm69znooKebv
yogm0Sa9h4GMq195YwJtiNMhkZz2RNbOtgwPIO+diBwuNd35J2Vzl3G5JMUTH+U5A/Asc1GeX2qdGxtDvC51vYf9ct8TqcPzMD4sWZke2/kwLYIvgUlACVkSTGl+aFUx
VlPpPG3ZuskyMvx562KhB6BTe4B3k/mbHjIUfqo67SIfXy7KnTBGEk0rgXVj2MzAi+klPv1jQYrqJD5P1flDBI4h3ubz/4TnDM0KGuQDTV7pwsN+Z5gRZVNc2Eu21Tpg
Ms6Yp83sbEijSPVFltsRMJ0Wl9N2kOxJrtSzwsuUoTweB5119q7F4OroEo8GyVII/fVihEy496AqRRQztv+S8WFSpK8LoSM34kzUGWh7HEThNQIwxRNfNJ5YfE+6CdJG
T0AdSo0+Ioxd3pOapgecMcqLgu9BiGogLtqZQaXzcU/iEj3iAcJWSeyJGc0PKR6B3sT/zw2Git/Qg3Mf8CMddKfX8jghJY2KiMFhN+T/UkwRqLQhyN1uhVIRyPITULae
nkPELMSQBI3KYVRngPExRiuZCpxaHbZZROUajL1cybsOhSEvMncJOxvvLDSGvNM88lW1k7K67w8sZ7RTf4mI5tmo+cwJby5CHG07RCJjR5zKiCbRJr2HgYyrX3ljAm2I
0vZ/C5D4uxV8hGR06yAxc9JXdM5YJxOsLcbMZcdwbiZmP0Vl41UBWqZtS2xqu2bBTQgpui1kSkD09TMlH3otg94LwyiXoYmarE4ZhOwZLlbLi9v4QNDxqu+7C6en51xj
2R3IH+x37LJn2vgK6C8A5mgpVbJCjr4V3OpcS2pe8oZtmhmbSQFu/4QZ3IQgMYQ4y4ucOVJdP1qgObTAZcYBa42sXL57daIMNSAk+4T0c8L14CGxtily+5U+nzoiY8iq
JAPf/bz5bE9s1ZLe5FFY2ChIBgLAU7dY0eVcZA2CNtH7rBWUj/jIHLnGrXXjRi/hQFjvGImy0+d2OsFkG1Ek70xPqKS5trQKu+v2WMqqZz72uzAflGXdSR4nP5/retPv
AdLXJI+tSBwBC+y44miZhrqOWVaXblj/fBFugf3xdf8zTHwCfWRG408mCWP0CV5TemTS4ew385msdNaYOxgOWcqIJtEmvYeBjKtfeWMCbYimMbKf63HLR5k+1IhTQZHc
elTZo7rJ6+FY/a9ecaejieP2FZREnRjNztP9isGe+bCYZzfYHTkVllCzG87DfQon2nwprEjEJ/BEkk9longSKYNxF05+fMMIhjTy+zEu7XtZEcVzu+UBm8LkDotdeQg8
tCEMWIDx5dms2kujiRYwRYa4quT8236u5UxHPnoh99xtvhBy+3cldQYYnzBoJ9eBXIA6IN7aK96lFqPI7XaeZomvX5jRYBoyP+S0/fQvdRrWVhbKmdFC/mAJZhygu5/R
d8j3axqQaW8FTnWHHmHrRmlsD1sr5eL3wxTUd1iaL0O53eHof1FA4ugep5cYeOtfVMaUMndBwF+kwMksXvheRkusv8CSPjuliVbdn4mYBCPoiyOgkzMOt0oYdBsF9wQQ
e3IlTH6FpMBuoPPAYFdjx6iupd0oW5VljSHWixzzLlKdYWHV3b4pRbC1p739SHkKcgcuqXz8VKFxDjVJUfNjdo88h+l6GH+gqgzjbxF3YXy/mR3czZGu62PbkK/VONVo
hMhbM9s0YrP3aHIgmqJs/XltsZewUmAVwgnxzRy9gYIuYpGIjaUi7tf3s84xauPrgRrInBgZD19HN9j5BZzno7yimkA62k89jNSABxu1GQOOXenBtQMYYzDihO2Ri12T
g+2eVqtBGxjRGZgyjSEzN8cEh43PVtce34eyDecmZXD7rICpy6vrQuFpgCGDT3b1682C0XI602dtdzg0zQpee8CrUx8bu5riiaYO4t7b5ThFWvHmKKf63yQJocUab9xY
HXFUaBdcPqFXsErURCkDjEj1C1wYfDJJ/EwGUKiy3SzTIZGc9kTWzrYMDyDvnYgcLjXd+Sdlc5dxuSTFEx/lOZ7CFBX0buYty3IPfnEQN2ztvIx0hi3glojzv68uM6k2
zUBH0P+b2ClmLFB+Gv9Cs4CyJiheCy37mgu1JC2h0Wnjp/+fY/tDq+DTCPeRLVk0H18uyp0wRhJNK4F1Y9jMwAwbOMQPYtpSfzu+EPqBo5JsWPwjGl7Evf/FkU4Os07/
6tV0ffa1VXNfoL+iRFGzU2vl5rihtV1SfJMjTund6wWUsmHTSZhXM5+/iAOPU4mAcdOwFk9lnsWLsL3/muCqVAPfZsPGWV65rUBDozqCMorILWZQpoWgA32jr9HoBvFi
GW4IzuNIWxMYqiD/fsRVK09AHUqNPiKMXd6TmqYHnDEDo+ZzUHRMyXKj3Q4IH7NqYeGfSHQJLgVLVA7s0K0WmEDbhtWBdAzEGqD4uoGyp3KTjc8duKCrlNNDZrxv2rrn
cjveAzO+/7U58YwS7JUaF55DxCzEkASNymFUZ4DxMUYrmQqcWh22WUTlGoy9XMm775ZaBlBLUuNVfn47ChEDAXkPLRXUou+liMJBuf7hZ/fKfrMjWWEGT23GKa8rrT/F
F4Ne3/tBSdh60ctPP9vbNapdTQe1P54xVOX2gkGNl9dYUV6xgeS0bEdikSLq3qj0n5RMGB2cEMCirr9o6qVWDs8oxwxhq9Ib5mKIG72IP9sCpVjkRPg/UslpcFUR5145
y4vb+EDQ8arvuwunp+dcY0Qirb4rkiYrRjK1lWYQVG9aLmnzDcx88l9Kw5LVj8RmbZoZm0kBbv+EGdyEIDGEOOcJlKqswZEEr9EBm4DjqjcNksduRJB0rcnFyMUed+9x
NmWWg12F12lg4BpNV1U8xyQD3/28+WxPbNWS3uRRWNjTzM50LafcyBCGavC0qamXs2ZHalXWLcl7vvP7DTzkEt6OOxecMHlXVdulD1ESI5VUnYDYG99HjGn10FyEDSBc
QMmqsJAIM6uAKSZME0akDNQuFzWpJAqAosAENCAkl6oESZq9HN2P82ntD0UYKmbv38oEg7oGprJ3iYpyga3KjgBYs0OWmRE+zk3EhghYWrnafCmsSMQn8ESST2WieBIp
pjGyn+txy0eZPtSIU0GR3DoLXOjJ6bdcpkMb7pacHt2s1fzkqRXBLlGUJWaBUgLeewzjflE8ccuOrTjfR5PMZvprREx5PlAIIKsuqCeWD4+DcRdOfnzDCIY08vsxLu17
++0Ym9qzeUUGTDAClc8vNEJDT8DXEZPV9GRP6vRyvefZUTx4uWvjRu0VRZMaHMl08PUZrvwHxt2PNViA2nWv2q6yZlCrv6VDhCYyIB1b83YAUFsO+IueluMlUWAiGDvP
RxH58+xPEcmMICwEfFs6D+GpxkTbzEHsDlCqC9zHU1SeIn3zbVuXdULmi+GItz77yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhLrL/Akj47pYlW3Z+JmAQj
EstAFfTRAYUadRdd5m7UFCcXTmjuZYedDF5Zh2NFM4NJb00XoIoG4ct2t9nx0Sr2CBFKc3zHy16oEUEMNaH3TXoptMq4JUw7PIguhdGP71aPPIfpehh/oKoM428Rd2F8
+3O/rJMij7UQnXoERuxubITIWzPbNGKz92hyIJqibP3Ujtq8y2CvINBje8YenfasCryAIMpuaGv58oKmH2qc9oEayJwYGQ9fRzfY+QWc56PC6N2gewbeb1w6Jweas1zk
pLdrasGdUNTAEhszu1+wQbabV2cNGISQcP+KupZ201OfHXC/bRo475erqvIc+MXI0vjyatqlCOINRHPb7mRDpedSvAVOygiBifDXV9Td56PssG8EJwvJW1buRvFagoBy
C4SxuoR0Q7n8h+pECBGYr+ciDPTnZZazCr2nLu1ibwui60aYd/LdYG7DxwJza9Cd4nGU1gXusKfbj8z5/LZobS413fknZXOXcbkkxRMf5TmDIVx1ZNlJAAZROJr0b39G
2xKVbWglVvs/Qum5AlqAtmDpvb7r68q35y41tG5ECgBeeUgLiTsuf1joWvvuJEVRoFN7gHeT+ZseMhR+qjrtIh9fLsqdMEYSTSuBdWPYzMCFumaGQBLvSsPkdP+XgSZ1
D0aW5ArJPqq4Q3ic8Byhomx74GoJyO9XEjmz77yLuOEY+lgkPoNPRKsGR3TFQ86lnRaX03aQ7Emu1LPCy5ShPH5dZffqmvlIgiIJ7o4vXPiYEM2mQJCY2V1bvVt/mz1V
RK6q0VoLiyzL4hM5mmYYx/Sx6xCahDz/qYe7Ju60j29kOsOEaslOzq27a855ePp0youC70GIaiAu2plBpfNxT0Lq/wrJM6YJqI8nHbnfcC1A24bVgXQMxBqg+LqBsqdy
i/7P8e7ESyfLyrpYbp24Yj06/CLwLe0/X9/NtTeJBlQnsol2e8FnsP6FJWBuVwVwK5kKnFodtllE5RqMvVzJuwqvCP5j/s3s1KpnGFIttb8QMRKs+M89biQvL/E3g/7W
UwZqFrmctMiWvohlxEGfRX8A/j75oRxgM/gBLozR09rS9n8LkPi7FXyEZHTrIDFzcLnlKWiJJ0YCwvzrkYFatTMYf6usFFsN3IHcbjqPoqJTpuA7aHOlUzvSIMDFGxtb
g2khQuDSakuK0bhPq/EA2j1u4jaleNdZJgOKoVARy5vZHcgf7Hfssmfa+AroLwDmpLU+d2v95+WB3zr9qrEGtm2aGZtJAW7/hBnchCAxhDjnCZSqrMGRBK/RAZuA46o3
g4PYD269w03GSQ2xSe7HRDZlloNdhddpYOAaTVdVPMckA9/9vPlsT2zVkt7kUVjYIeyc+CGFGIT/xuT+zGXc3T4hCguqiTViQ+TmdiVlEECOuIRRooJs0sb997/120mV
rfYKQiEK8VpsOKtzmt7ze/a7MB+UZd1JHic/n+t60++gW74SqiykSlecXd4aSeGA3bnLi12y8qwu94R31X8OmN/KBIO6Bqayd4mKcoGtyo6t7CxhCOwT3raYRg5LriTq
mr4MnTQzL8u5Cq3DgpmjiaYxsp/rcctHmT7UiFNBkdx390ssHHW9bT9EqbhChWA75CJxF58DwuP+KzXN5XTAw6w4HGns5yTPlrVLa51nHdyMIh2A0TjlVhNEnan2OChw
g3EXTn58wwiGNPL7MS7te1kRxXO75QGbwuQOi115CDwYBeaDGR/7u9ZXunq17CGvhriq5Pzbfq7lTEc+eiH33HdYgplxnjKBcpmuMnAqwa/afCmsSMQn8ESST2WieBIp
ia9fmNFgGjI/5LT99C91GkcR+fPsTxHJjCAsBHxbOg+lfKDVIJ9rJfeW/irISIK0IYwZoQb7rLTDvzin/7ZiC5L5oQj7lUrrZ0XKnjXlSOtw70Un1Q9IUc6G91GseXXA
S6y/wJI+O6WJVt2fiZgEI1IGASDXJ+j/e7SpF6VUXtOGmi80V9ocuwEK8kyA+4Nrs4+auKDpDRaaAlDwlnNoYm9YfP+hng+lycaD1fvQWMhkJKoHC3IKer9WUkT3GW4B
erZqgp/njJBc4V9mdMoKON4c4SxbIuFKqFpAzkUkZD6D/qIOKbPGmxLrYvPhdKMcWThhSoxDjYNybNuJtXmYkAcHf763heL9QB1pkvJazSpVEEC5mMRS920Zx8nelqEy
wujdoHsG3m9cOicHmrNc5CHvIzUVnQj5Ql0vw0Kkgh2D7Z5Wq0EbGNEZmDKNITM3dZoEs0u4NqWaBdbD6ClOevusgKnLq+tC4WmAIYNPdvXrzYLRcjrTZ213ODTNCl57
lW1MPrFtyZUbU9Jcprku6EVa8eYop/rfJAmhxRpv3FjnIgz052WWswq9py7tYm8Ltuj/CtKPJY6G22YjImQl+cnAnk/AkTdsC1rlckf9aSkuNd35J2Vzl3G5JMUTH+U5
y79FSrvtO/zhxn6tr7yDqNsSlW1oJVb7P0LpuQJagLZxrEJWOMNee2yilas7avaW5XZ9MWODE5yfGrzxiy+zfOnHVftzjYQ56eym/QM73EIfXy7KnTBGEk0rgXVj2MzA
XxgFerwuOSqgdwURKgNy6mxY/CMaXsS9/8WRTg6zTv/gHiLOYBsmnpvuSXn70ruGUitjiYWfbCE9/vBr8/8b5JSyYdNJmFczn7+IA49TiYBq1qS5XiZzoeSX2s7UPYlR
wzL73tawU1fcJnkuZ9rwF8gtZlCmhaADfaOv0egG8WLVpehx0zpgot/QYNZtc+jvfI8M0R3KqGr6cHMXtkSzeQOj5nNQdEzJcqPdDggfs2oxThnmr2jYVz56qGorr52Q
QNuG1YF0DMQaoPi6gbKncjZDEASYRD9NbEgYG6JmCtwMtRQW/5bjYEzz8yMKcL95oY4ZFtMWUeI69RCmMkyCzZtxm6kiQNLA4JcB93Vx0eTafCmsSMQn8ESST2WieBIp
eQ8tFdSi76WIwkG5/uFn99t5Xw56sYXOIK0XKEHYHAzKiCbRJr2HgYyrX3ljAm2Iql1NB7U/njFU5faCQY2X16AA7z0uCCwY9P3VVS5s21HfVvMNN4aFZPRb6ILq+974
qC8FN8TpnE/kVLIpmNKkJTVfU1Ef2zESal2+E3929yJ8aTcT+LAmjL5Mqt6/pmdN3A/HQUAYHGYwc9euKnMf/G72B0zJbtNS/KendGthYGxtmhmbSQFu/4QZ3IQgMYQ4
3gviT5Rm++4A+a/sW24LlxHgu5D5rCjEGSrALpqJYvc2ZZaDXYXXaWDgGk1XVTzH4uI7XurWdxkjeOumOwPlbYXvEs6ey6FxshFjuObyhyKzZkdqVdYtyXu+8/sNPOQS
b5YqCa3uEhIOLnyf3uDDtTLOmKfN7GxIo0j1RZbbETBAyaqwkAgzq4ApJkwTRqQM08p7TTPLBqJZNeriWVcpHHHppJYjgpGkgXvbawejv+9JgAJITpEM0ere2AIXGJJL
FLj8lY4TmE5Twmk7VB8YalTGlDJ3QcBfpMDJLF74XkZuE8JomAdCaF3g9Zf84UgZkDpXiWvVYbYIvCi/TnfMh+QicRefA8Lj/is1zeV0wMONDF7MsCzx9YzLKRytBIB3
TgT4QtMKn2r4tAPdeNFPfoNxF05+fMMIhjTy+zEu7Xt+l20od+UaDo0ko4eGEnF/zNWmJC9UOX95bjk7NVeePYa4quT8236u5UxHPnoh99wvaoRak294sEnpfRKH1KWa
/TTrXmCv0PNeRPJn/u1LbImvX5jRYBoyP+S0/fQvdRrJs89YaScMlSW/2lahJdrjz02asvNXIcjRDnE6QiDYMjDacDRbVRBi/68EYfSvcaPvEqdk4LOonqk0MOhy/7Ar
VMaUMndBwF+kwMksXvheRhJGqJWn1t/qGroimMFAGFYsocFuCt+Kg//Fm74sEUE8juJDucFoqH6IPHRppeAeAORoNEyh5SiDzX48QX8wWSUiTiOve2+wgxyxFcmEqMkZ
cgcuqXz8VKFxDjVJUfNjdgYBZKGW20y0NuyBLre4D5EoWOauwIEEtTEb2Xa0cPovhMhbM9s0YrP3aHIgmqJs/VOfhWCOswRDbSrPx63rzDEwpL2qOvwOFuI/3x7cQf5K
fUgoSjZJ0mfLOvTfraoVzkFbd6TtX/uFoAG40CPc9JjPq6mvdB3NU8ftvbYWcxNjCv2hKWXn/scQqFxHS8LBCJpbEdA2xsIcQBfgFbhYA5NuPcqjj4KMfzKD264bGZmd
HnxxE58x7qzsr23/eeD5ypXjcPCNWLHj8MyKWXpjaEDw7haRU2FIPEVTdfREZzeLVdmgwS2YE7P6+awFzsnabw/OGG7gfoM2xpCtShQnGsbTIZGc9kTWzrYMDyDvnYgc
kjcNPXBp4PFAtM7mq3J81X8A/j75oRxgM/gBLozR09rbEpVtaCVW+z9C6bkCWoC2xLtr2qEIGqj24LUgJ2uxsdzB98jR0TzjJrgFdyQttTPpx1X7c42EOenspv0DO9xC
6YI0BiF/vUm2oVbBPuUF6FMaEHlsnQsQyKZVFILUEq9sWPwjGl7Evf/FkU4Os07//NpjZMHdA5MRgX4htPt3vcqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqh
g3PXt6rrm8wh6BIuwAsZ6lUQEhoK217dO6xwx3++2wksX+bKTugLpOfqbyjby6quyogm0Sa9h4GMq195YwJtiE9AHUqNPiKMXd6TmqYHnDF5l4tHAQTcyKdVO4u+Yagg
4/cZD5qaXN6DhKB+PiGL1UDbhtWBdAzEGqD4uoGyp3KcUYiALcUcFefnb8w4/SP4LnfpZMUMik0jsG/ygpO4HaGOGRbTFlHiOvUQpjJMgs3QPqm7LzmyJiimOGB4VGSF
gC8/AkNK4iytXUzIponOA3kPLRXUou+liMJBuf7hZ/fS0n/p/9Gh992n1gn0OvZJMs6Yp83sbEijSPVFltsRMKpdTQe1P54xVOX2gkGNl9eZuusOS+fSEmY1PeniY/fE
SZXdRwN4saED/s81w/rdTKgvBTfE6ZxP5FSyKZjSpCUDmmGBJczo7pl5Py7I9xK73gRHoQ0bubQUMPVuAEVMOitPQgGgvhnT6E6HCAMb+XhHhCTV5kDXCeZNfRIkkCQ8
bZoZm0kBbv+EGdyEIDGEOEbKLGLn8rBnOqQ5+REJJtAEaJJLqbX4XZkB4zET0nRp9eAhsbYpcvuVPp86ImPIqpG4hFclJcRLbxcCqfx48y9w70Un1Q9IUc6G91GseXXA
s2ZHalXWLcl7vvP7DTzkElPf9zXccrZsteeLLUgMz9fKiCbRJr2HgYyrX3ljAm2IQMmqsJAIM6uAKSZME0akDLyPVXrCdZE3VELCpDEucLkc+TaNxDDi/A0Bd7t7rbQA
O7sI1CYfGv5Qb4MUHSCxkhk8USwkW34n+ns1trJ9OWNuPcqjj4KMfzKD264bGZmdRU7c4+AcsoCp8kKEqxqyMkjGwpX1xVupz3pPEAag3QhHslolreVfipthc+zo1Ki5
d1/dbi1L2ORRcwHXjV4fhGt3+HddpNoLrTwrdq4Aa/yDcRdOfnzDCIY08vsxLu17UJDn9h522Q4n5otk1oHXodp8KaxIxCfwRJJPZaJ4EikvKAjSdz+er6sZXFxlkQmb
THNI5UIdnGgUA28z3bNMxMqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13LmRsA1d3SBGos7+fAsg0FHNiMYD8eF9P3gXRMPHskkYgw2nA0W1UQYv+vBGH0r3Gj
aOCfoHtDORRG/pGrbsssQMqIJtEmvYeBjKtfeWMCbYgSRqiVp9bf6hq6IpjBQBhWDrF2IMnl7VSYWTBbnGpI1o7iQ7nBaKh+iDx0aaXgHgDDdKiRPeZLGHR5xVUPi7Si
vwY7sko24S0fR0QZdkCxenIHLql8/FShcQ41SVHzY3bMlrA6kAKGmalSZre6myAHQlS7ZlihHgCaTRamVg3WgITIWzPbNGKz92hyIJqibP1LTdOUWjfxjuucZkifSHJ5
yogm0Sa9h4GMq195YwJtiIEayJwYGQ9fRzfY+QWc56MqozDo2RCt9t3uNpPiDHMswrrP0/aYg3mgzNjm3wiXCSzhwJRvtZp5VVnKhTjqk28wXz7HPDGZeL/rbKK605AV
yogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh0aiuEUqiGXSR48Ux4POgj98O4WkVNhSDxFU3X0RGc3i5LKQpkDwkcQf8KlG6wH9eouYpGIjaUi7tf3s84xauPr
0yGRnPZE1s62DA8g752IHOwgBk7QhAilwQTBAKROVLNNrOe0POlmnvEHzG3DuAc+7JukIBvhL6aNiYGSTNKtvE2s57Q86Wae8QfMbcO4Bz7KiCbRJr2HgYyrX3ljAm2I
oFN7gHeT+ZseMhR+qjrtIoU2knnEs5OCk04qUddxYB8uYpGIjaUi7tf3s84xauPrewRCIRmd9fsmH288aAUGOi5ikYiNpSLu1/ezzjFq4+vKiCbRJr2HgYyrX3ljAm2I
D7YfOYh4V9obUTgnsMT8MXUAnUCmR0X+/xWoUE9QxtFdociG51a3adP6dskgTld+UAyR+GstxIGIgFg/xIL3qUEeEMhggIZX1RtHECuZZjsFTNf+juK880vz8jdPp0Nw
ZeRVCx/7rQkiPMyXxzciX8qIJtEmvYeBjKtfeWMCbYjTIZGc9kTWzrYMDyDvnYgc80s1u2OqHYTm0Fd/2Mp/6N4dUnit9vxzk7l/HYQFUOmEyFsz2zRis/dociCaomz9
4AgNDv3zl0QV75nL2CAdEbq7rpYcmgzHjQxFsY6vd37KiCbRJr2HgYyrX3ljAm2IQMmqsJAIM6uAKSZME0akDNRn1JQPcRZihGp83Flix21Jld1HA3ixoQP+zzXD+t1M
BUzX/o7ivPNL8/I3T6dDcMWJTIIcCr9LCwa/NQc13ZpUxpQyd0HAX6TAySxe+F5G0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+gRMOuCN8h1grwpr/xigFit
LdevBXBm+elemUyDJUCVKL/k52cysYmRiqukdE1JEf+W8MwpU8uF2Z3WqQjTVPjzyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60++zbCGM04VIKW7e+SwNVwIH
4z5DaZW/k+0+VPqbqK8s3QVM1/6O4rzzS/PyN0+nQ3AviTi7UulykOBlj2eO2DgdMs6Yp83sbEijSPVFltsRMNMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o
2EBgpX/NKy+lKfUNg+koby3XrwVwZvnpXplMgyVAlSi/5OdnMrGJkYqrpHRNSRH/SW8tEgNwizg/aIHPmsTwucqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
l0tZCyTD4gdmV6ID04hR60mV3UcDeLGhA/7PNcP63UwFTNf+juK880vz8jdPp0Nwxf0Ji4ClVM7OV2STMIRiam49yqOPgox/MoPbrhsZmZ3TIZGc9kTWzrYMDyDvnYgc
80s1u2OqHYTm0Fd/2Mp/6LT56Es9m4ebg0VXf+fiydot168FcGb56V6ZTIMlQJUov+TnZzKxiZGKq6R0TUkR/7uRkxvR8jmt/P/uHxXrTJXKiCbRJr2HgYyrX3ljAm2I
9rswH5Rl3UkeJz+f63rT72fTVfpSEbDI7UItikJJantJld1HA3ixoQP+zzXD+t1MBUzX/o7ivPNL8/I3T6dDcJSolraezAT8nrNfuhCfocrKiCbRJr2HgYyrX3ljAm2I
0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+i2Z1Pn9pz9CCDpAxSYE33TLdevBXBm+elemUyDJUCVKL/k52cysYmRiqukdE1JEf+Z8nEW9Kwu+bz9vsluAFdM
yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+/tx+B7hL4We6zxndKWymIDSZXdRwN4saED/s81w/rdTAVM1/6O4rzzS/PyN0+nQ3DrmJEJte+kgqmNkbMG0gbL
yogm0Sa9h4GMq195YwJtiNMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/oMYn48LU0q1T0DwkEVyp7jS3XrwVwZvnpXplMgyVAlSi/5OdnMrGJkYqrpHRNSRH/
tiqPF3ZUmtgfqH76MQqRJMqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPvaKwy/vLcSjXTbtgS9z3te0mV3UcDeLGhA/7PNcP63Uy7MLb0XC9WUirLL562h0f8
CRBl9MQwBik9LJVwV7C1AYtga29j9WzWHanK0tEH3sTTIZGc9kTWzrYMDyDvnYgc80s1u2OqHYTm0Fd/2Mp/6DAjKrP79fbP6Ik2gMlU49uEyFsz2zRis/dociCaomz9
4AgNDv3zl0QV75nL2CAdEemljNpSaMX4LB5WwQ3hGOrKiCbRJr2HgYyrX3ljAm2IQMmqsJAIM6uAKSZME0akDJburv94oVHUzXiljpsJgAtJld1HA3ixoQP+zzXD+t1M
uzC29FwvVlIqyy+etodH/GZovmyHAqJS/dqDd4iuSMunHqOgU55uXDWCN1Ydicbs0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+hD+Qd00v/wS6qAzebfDDpZ
LdevBXBm+elemUyDJUCVKJi9qGIlLSG/uFN5+JjTifEQXk1WaztjxA0X6rG+lJ3Ayogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+/yyL0Ob40/nxXitw7Q/aeC
SZXdRwN4saED/s81w/rdTLswtvRcL1ZSKssvnraHR/yaHfoX+5a2LrFlw+wsYIhoQSZpSFO2o1eAup2K2DYwl9MhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o
jl3pwbUDGGMw4oTtkYtdk4TIWzPbNGKz92hyIJqibP3gCA0O/fOXRBXvmcvYIB0RhApa6QAxR9CQUDD4YFCYsMqIJtEmvYeBjKtfeWMCbYhAyaqwkAgzq4ApJkwTRqQM
gpNSX5tPo9YFbWFvZI6XTUmV3UcDeLGhA/7PNcP63UzFpwmvhH1+C9P78UWLfY5Yyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjTIZGc9kTWzrYMDyDvnYgc
80s1u2OqHYTm0Fd/2Mp/6KJHw7fK7CTEw1FQq0fJvvWEyFsz2zRis/dociCaomz94AgNDv3zl0QV75nL2CAdEUZPCECFOonJJOpocqHgW64mZ9Bzkwz5KZShD3A+7aLp
QMmqsJAIM6uAKSZME0akDJH9wEzooq+fUsQw3xpXFphslZJ6MC1ETrwwkJ/F7F0gU6bgO2hzpVM70iDAxRsbWz2UHhRP5OuAUuUz9JhC5sAHB3++t4Xi/UAdaZLyWs0q
HA2EDF+ychpMfvoMbyhrOP0NwjVoPQpcuqk5KJIg11iK9iSqp1HId/Prb/+GduBMLdevBXBm+elemUyDJUCVKKudKnSHFFnogOY+sKZafFrd93Jg0pPUijZXofrfCAqh
yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+9sOgrzMFFK9909MbNiwRQD31bzDTeGhWT0W+iC6vve+FOm4Dtoc6VTO9IgwMUbG1s9lB4UT+TrgFLlM/SYQubA
VOF9g7sh94P6znjjyr4gqtMhkZz2RNbOtgwPIO+diBz9DcI1aD0KXLqpOSiSINdYU5ik5dVm1fmlp1owVld8Vy3XrwVwZvnpXplMgyVAlSirnSp0hxRZ6IDmPrCmWnxa
z8zWxJy0VvLqpsRitwmtq8qIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPvJee6+UvDm8dKHT970fcGh0mV3UcDeLGhA/7PNcP63UyaMuBAGBEB2xeOGnMSsijz
IG/wGYVQlx9Uz/bopuLEb8qIJtEmvYeBjKtfeWMCbYjTIZGc9kTWzrYMDyDvnYgc80s1u2OqHYTm0Fd/2Mp/6HbX6W1L2UArFj6ZjZvCgYQt168FcGb56V6ZTIMlQJUo
q50qdIcUWeiA5j6wplp8WlZT6Txt2brJMjL8eetioQfKiCbRJr2HgYyrX3ljAm2I9rswH5Rl3UkeJz+f63rT7+V7j0Mvob3xonJhdB7kyqFJld1HA3ixoQP+zzXD+t1M
mjLgQBgRAdsXjhpzErIo89UZX9LXDIf0n/etQsgSwWLKiCbRJr2HgYyrX3ljAm2I0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+gy51IgcF6/b2UlxZUevH/c
LdevBXBm+elemUyDJUCVKKudKnSHFFnogOY+sKZafFrAgkmPjGDrWZ9z3bg+iKrSyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+8dk+RqpSK5bqK4BPCi5LXz
Am5HG//yPBtVhcrExLB3xJoy4EAYEQHbF44acxKyKPPSX2Oz4H90SNdFRkyKUUrxVMaUMndBwF+kwMksXvheRtMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o
foYJ4iG+s5GBAS4gdC+Ngi3XrwVwZvnpXplMgyVAlSirnSp0hxRZ6IDmPrCmWnxaoUTeXg/41jGKjYKdkBB6LsqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
rxwRGkx0NXMhr3apDSRa0mOmZu33Oc9RgiStST47G/maMuBAGBEB2xeOGnMSsijzgnhMia4omX8FtxOiEJkaXVTGlDJ3QcBfpMDJLF74XkbTIZGc9kTWzrYMDyDvnYgc
80s1u2OqHYTm0Fd/2Mp/6K6tve0DFPWXXGGJmVLbYN0t168FcGb56V6ZTIMlQJUoq50qdIcUWeiA5j6wplp8Wv2WDCF+p5mlC9wYGpid/33KiCbRJr2HgYyrX3ljAm2I
9rswH5Rl3UkeJz+f63rT7yNYaItfH8R6Y0XbnxFRhiJJld1HA3ixoQP+zzXD+t1MmjLgQBgRAdsXjhpzErIo82kAQwtzExifETAH71bpkrluPcqjj4KMfzKD264bGZmd
0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+gh7yM1FZ0I+UJdL8NCpIIdhMhbM9s0YrP3aHIgmqJs/eAIDQ7985dEFe+Zy9ggHRFYLPWSx6pzGKmi2XjFgJCi
yogm0Sa9h4GMq195YwJtiEDJqrCQCDOrgCkmTBNGpAxQuxrj8/lZp/iVWaiHCRc5SZXdRwN4saED/s81w/rdTBJQ3HewjrZ38uwFP5ZO5s/KiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiNMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o6FUFXDi4YxAGl5DqmzmcpoTIWzPbNGKz92hyIJqibP3gCA0O/fOXRBXvmcvYIB0R
zGt/K++s6vlPaxt8YURdvWOLKN/NVM9esVtn30j64slAyaqwkAgzq4ApJkwTRqQMDYbWiAHm20JylrdbPLbJFEmV3UcDeLGhA/7PNcP63UxTpuA7aHOlUzvSIMDFGxtb
PZQeFE/k64BS5TP0mELmwGWRVbqy/1te0y6uDxS8QBjTIZGc9kTWzrYMDyDvnYgc/Q3CNWg9Cly6qTkokiDXWMluNWh6NU33fn0l+muMJeiEyFsz2zRis/dociCaomz9
4AgNDv3zl0QV75nL2CAdEVKreb1Qn0kFSmpGwZFI3uIyzpinzexsSKNI9UWW2xEwQMmqsJAIM6uAKSZME0akDLJfeFOaQbknyYPAh4IEeSxJld1HA3ixoQP+zzXD+t1M
U6bgO2hzpVM70iDAxRsbWz2UHhRP5OuAUuUz9JhC5sAzpu9l3dXPx7c1mv75CSFs0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNX2/xiQ9k8L/ABz6nNLGSu2
hMhbM9s0YrP3aHIgmqJs/eAIDQ7985dEFe+Zy9ggHRFjZjk0Kw1F1vQ35yKbepTNyogm0Sa9h4GMq195YwJtiEDJqrCQCDOrgCkmTBNGpAzbzLrrhf+tRr/73LF7yLyX
31bzDTeGhWT0W+iC6vve+FOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLnD7E/9kne4PLvL/kIw3RZNtMhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbg
AfJJVAe02upn+P4DNeQ7lITIWzPbNGKz92hyIJqibP3gCA0O/fOXRBXvmcvYIB0RSsRu0eRvjRWI3hXEj5Jtq5ZicKksc3MYALhdLrZ+0R5AyaqwkAgzq4ApJkwTRqQM
JuWqsNVvk6tfHHQCDTQpF0mV3UcDeLGhA/7PNcP63UxTpuA7aHOlUzvSIMDFGxtboyK6GOi+0Of+omugCmqf+IcLT1BKq6WHmmjLJ5Ew6OzTIZGc9kTWzrYMDyDvnYgc
kjcNPXBp4PFAtM7mq3J81a3QjooRma47KJl4X4OksTCEyFsz2zRis/dociCaomz94AgNDv3zl0QV75nL2CAdEf8ia2ms1kTrKqdxmywLJ3IIHI89GHO7Fgaiqszij2Yw
QMmqsJAIM6uAKSZME0akDNWkEBvZJwHeE0p0KZnL3zRJld1HA3ixoQP+zzXD+t1MU6bgO2hzpVM70iDAxRsbW6MiuhjovtDn/qJroApqn/itywArBa6dMsMhQctS6nCg
0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNVs48gRpjUSMHwljLGeSnDRhMhbM9s0YrP3aHIgmqJs/eAIDQ7985dEFe+Zy9ggHRH4rOiksy05VcGdaqk4UZCh
2JSh+UKRKMPsKIdv5SksJkDJqrCQCDOrgCkmTBNGpAwq5GCz/pxxirrLTSaKVFGBAm5HG//yPBtVhcrExLB3xFOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4
H3Cpn8ft2iEQ+fEAfKIpbtMhkZz2RNbOtgwPIO+diBySNw09cGng8UC0zuarcnzVimEhNhFMkiHDLrUSaWCDx4TIWzPbNGKz92hyIJqibP3gCA0O/fOXRBXvmcvYIB0R
kLi8vTMYGfOsgRqwF/sSOMqIJtEmvYeBjKtfeWMCbYhAyaqwkAgzq4ApJkwTRqQM5Szz/o74T+/F0BNe27YxjGOmZu33Oc9RgiStST47G/lTpuA7aHOlUzvSIMDFGxtb
oyK6GOi+0Of+omugCmqf+NlS1V0pg16vtF17VbhT7sbTIZGc9kTWzrYMDyDvnYgckjcNPXBp4PFAtM7mq3J81U3+C7F5PVEBnmRkBlnc6qKEyFsz2zRis/dociCaomz9
4AgNDv3zl0QV75nL2CAdEeP5B75XmukM5kAVkovrdh4yzpinzexsSKNI9UWW2xEwQMmqsJAIM6uAKSZME0akDP3Gk27g8XFocmIEhA2rsrpJld1HA3ixoQP+zzXD+t1M
U6bgO2hzpVM70iDAxRsbW6MiuhjovtDn/qJroApqn/g/wL09aUNgISFLweRcjRav0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNWelWAGd8ZpgT5HRsec5BNx
hMhbM9s0YrP3aHIgmqJs/eAIDQ7985dEFe+Zy9ggHREi2EpQUtX+XzFUyQfBsDb/yogm0Sa9h4GMq195YwJtiEDJqrCQCDOrgCkmTBNGpAzgA2osp0/mQ5OAA5D/vFDj
SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLn9E34thKlpTPJMUEB+u8QBNMhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbg
24WG0h6YlmtvZuVO1t0hooTIWzPbNGKz92hyIJqibP3gCA0O/fOXRBXvmcvYIB0R7NgRh2giE90bgrbs4VBhvmOLKN/NVM9esVtn30j64slAyaqwkAgzq4ApJkwTRqQM
bg2b5pn40Jpvfg7FRec+LEmV3UcDeLGhA/7PNcP63UxTpuA7aHOlUzvSIMDFGxtboyK6GOi+0Of+omugCmqf+EXTxpXDTFGmSVa05wJaGE/TIZGc9kTWzrYMDyDvnYgc
kjcNPXBp4PFAtM7mq3J81RjeYSm2VM34dabATX+7JjGEyFsz2zRis/dociCaomz94AgNDv3zl0QV75nL2CAdEav31grIlEvgec5EcJ2lZZfKiCbRJr2HgYyrX3ljAm2I
QMmqsJAIM6uAKSZME0akDEXcDHnRs4Qsg4X8YWp/afhJld1HA3ixoQP+zzXD+t1MU6bgO2hzpVM70iDAxRsbWxyLJM9m1+hZpHDVGPttMueJv6SaS85rhPoQfXA8fT6n
0yGRnPZE1s62DA8g752IHLnP5Pjl4sHgFuRC5wOFZuBI9QtcGHwySfxMBlCost0shMhbM9s0YrP3aHIgmqJs/eAIDQ7985dEFe+Zy9ggHRGY92AaxFzZItZdWL4Ux3Q3
yogm0Sa9h4GMq195YwJtiEDJqrCQCDOrgCkmTBNGpAy8j1V6wnWRN1RCwqQxLnC5bj2iK1Ds8eSRrYopgplH/VOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLn
iJ4o4hQdGJLjdN0bmtKjCpo4Ifv2lep3B+ga7ojdjKa5z+T45eLB4BbkQucDhWbgt/2/e7VsI/t6bVdgNw2LSITIWzPbNGKz92hyIJqibP01gPYvUAmz1OQefQ+Zb0QP
S21HZrlnuPkLTbU5mfuZAnLZMYECF1mr9d0WMpFXfPQ9/bEy/2EhLO01p8EQaqyAcBV1P+ORgIh9qfl5PT8eS0EeEMhggIZX1RtHECuZZjtTpuA7aHOlUzvSIMDFGxtb
oyK6GOi+0Of+omugCmqf+G/Pex2QFmAzaVGeGb8Wvu/TIZGc9kTWzrYMDyDvnYgckjcNPXBp4PFAtM7mq3J81Vw9sfeZjalSEPIi1hfaeCWEyFsz2zRis/dociCaomz9
NYD2L1AJs9TkHn0PmW9EDx+GpYR8ADrOY6tKpzL+3RCdmay6ovqVCrZGH5f9b5v19rswH5Rl3UkeJz+f63rT75pccraHocdEUizKU3A6pAZJld1HA3ixoQP+zzXD+t1M
U6bgO2hzpVM70iDAxRsbW6MiuhjovtDn/qJroApqn/iyK6p1kQ6EMqlBoI4+fj3x0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNVymm1mx9E8kkT27ky/Dai0
hMhbM9s0YrP3aHIgmqJs/eAIDQ7985dEFe+Zy9ggHREEw5o/kvPkuMCNNrmiPklcVMaUMndBwF+kwMksXvheRkDJqrCQCDOrgCkmTBNGpAyBPA1iqk8y9ICnDM2xMG5H
4z5DaZW/k+0+VPqbqK8s3VOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4CKPbDCz6Re2QgnqljnrfTdMhkZz2RNbOtgwPIO+diBySNw09cGng8UC0zuarcnzV
qdPX1/gYO+3Xs7vQRSyBJITIWzPbNGKz92hyIJqibP3gCA0O/fOXRBXvmcvYIB0Rvy4/uS1Anj1P+Mbj+aTjnTLOmKfN7GxIo0j1RZbbETBAyaqwkAgzq4ApJkwTRqQM
c0jR5ngpqUlcaRkgLEPU2kmV3UcDeLGhA/7PNcP63UxTpuA7aHOlUzvSIMDFGxtboyK6GOi+0Of+omugCmqf+LsSF2p81cOt5xXkVe3vpXfTIZGc9kTWzrYMDyDvnYgc
kjcNPXBp4PFAtM7mq3J81R4WIxwl5Gfyp+chdzZcCBSEyFsz2zRis/dociCaomz94AgNDv3zl0QV75nL2CAdEX+3zycJXv3XugBYn2Iq7j05bBHmYOQtmQPF0Dbqccjs
QMmqsJAIM6uAKSZME0akDGeSiPKbDL9LWRBPVx+U4nlJld1HA3ixoQP+zzXD+t1MU6bgO2hzpVM70iDAxRsbW6MiuhjovtDn/qJroApqn/gJ1PHrDtOquttelOkGpz+l
0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNVnYGrahSV2iRZiJA34nWcfhMhbM9s0YrP3aHIgmqJs/eAIDQ7985dEFe+Zy9ggHRGb/QEGak/JjOsKv3m77oBN
d46GCrXHO8eMAlHn80c6HEDJqrCQCDOrgCkmTBNGpAyghx1Fe59yaRR+Bu/Hfzl+SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4
ibHBEkAbo/d56M5JyNGQudMhkZz2RNbOtgwPIO+diBySNw09cGng8UC0zuarcnzVd22hlotPlSczGpCizzlbb4TIWzPbNGKz92hyIJqibP3gCA0O/fOXRBXvmcvYIB0R
WsnQVe1MGqIa1VMe8Dr/P9iUoflCkSjD7CiHb+UpLCZAyaqwkAgzq4ApJkwTRqQMg5J/pNvfVVYZA9wgCcS0C0mV3UcDeLGhA/7PNcP63UxTpuA7aHOlUzvSIMDFGxtb
HIskz2bX6FmkcNUY+20y56fXS8BvsWiMVotdhgWJS2zTIZGc9kTWzrYMDyDvnYgcuc/k+OXiweAW5ELnA4Vm4BJDKUj667mckBaCM6k2oMqEyFsz2zRis/dociCaomz9
4AgNDv3zl0QV75nL2CAdEYT0enC+em8umcqWs5uPjWTKiCbRJr2HgYyrX3ljAm2IQMmqsJAIM6uAKSZME0akDPewdiXoQsYOiNNUp80octhJld1HA3ixoQP+zzXD+t1M
U6bgO2hzpVM70iDAxRsbWxyLJM9m1+hZpHDVGPttMucIOamPWSJ/XpR70WcFHME/HA2EDF+ychpMfvoMbyhrOLnP5Pjl4sHgFuRC5wOFZuBQ8gJ62UO/Ww9e281lkRt7
hMhbM9s0YrP3aHIgmqJs/TWA9i9QCbPU5B59D5lvRA83urMCyR4nUKup2U/KBNU8ZXFcfBagwcC1Y3a2YDAWtva7MB+UZd1JHic/n+t60+/8UmSIfNhiZxzKAVWc1TKB
SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLn7Vp2xUlg7+JuHPKclm9kgCceyR8H1C6w6XaqOhjgzHa5z+T45eLB4BbkQucDhWbg
w/F+tWIMr5G7AYfvsYvpsITIWzPbNGKz92hyIJqibP01gPYvUAmz1OQefQ+Zb0QPN7qzAskeJ1CrqdlPygTVPNcnimzwEO0GEmyJ6R+6ZJL2uzAflGXdSR4nP5/retPv
ytSvGD4Z5Bg8DwwBsuMmtkmV3UcDeLGhA/7PNcP63Uzcg++/X9x/CCkPPmHMR5kEyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjTIZGc9kTWzrYMDyDvnYgc
zeIuhAoje7om6wQGQmm87Dm9Lc66zmvw3hphF8yJlBC4FhCnhAMb2C3XhmdoVfCtyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
9rswH5Rl3UkeJz+f63rT71HCbZN3AW36QloklgT2oTNJld1HA3ixoQP+zzXD+t1MFQgud5e0U76HRqctBOPJw8qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
0yGRnPZE1s62DA8g752IHLEuIFvwiCfdqBqGg0RLwUXP45sqZ4YalKRdnWUMnbqahMhbM9s0YrP3aHIgmqJs/QP81xEf/yCOtXCmcu1t9K7KiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiKuRCXjuaWzW1xmYO4DehHxZkzhIkNPb4bn2ZNh7cG0PuHHTshDjLlTcYXipsL37ajytD8f4KHDoyaK1cn3UWwJFLv5skCT5FvcKOqgzEtAj
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAy6UZZ1a+5OkLIbJ7LkepQHmXi0cBBNzIp1U7i75hqCDGv8jyfHPIiLSdovnsBzVm
FJqAD3lIDMFTIw5+HZUauYaLS7CveEpqs3M6kDDdad/KiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oUhd5pCsfLJBrk6auAEQsAD
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAnMZs04C9HXUfAVuhha+pcXmXi0cBBNzIp1U7i75hqCDX46mu0kAtU+cH3waQlT0D
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtA8irBFiq5/W4AZPCCvyETtXmXi0cBBNzIp1U7i75hqCBJ4uvjYoMWhumX3L2JyNV5
pZRe4QmM6mwnB4taJC3gHjgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAm4B3Ag2D3p4w7bSNc2ntyHmXi0cBBNzIp1U7i75hqCBSck51MxClvHJDPbACODmU
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAl3rLg6o85yqXYD++AAzpQHmXi0cBBNzIp1U7i75hqCBg2b6E9AN5aKoFxyw1wfU1
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAh7hVnOz5PUBHuu2BlW1+f3mXi0cBBNzIp1U7i75hqCAgXRcSWzE9RK7PoVeHSN89
JMu/mIob71FrLh75/bwN8jgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtApMLY1PcjjfSJ9uXb05pe5HmXi0cBBNzIp1U7i75hqCCJJ4o/Bh08A3eTSIRmDXHe
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAycyLZmANr31FpDWc84nQHHmXi0cBBNzIp1U7i75hqCAPmF0fI0JAB9RbwMPHyM05
1zV7SJMYIHpXwQ44MP2OgjgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAJ4xe4QlHxrcOE02p/Bz4vnmXi0cBBNzIp1U7i75hqCB7K6boorjbz4Tcw8dXbgW2
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAb2PYyGMm9wL+BfnRiHJFZnmXi0cBBNzIp1U7i75hqCAnq5Z5WkuquRpUo6KivdpX
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8F3d4K8YAznhqIv3pBl8DtAmaocPx8tshJHoaPL/9T313mXi0cBBNzIp1U7i75hqCD25wXoedIw4TvqHiiwDf+K
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAy6UZZ1a+5OkLIbJ7LkepQHmXi0cBBNzIp1U7i75hqCBBAFVbamuq6rsdaYU58IHl
FJqAD3lIDMFTIw5+HZUauR/+ImyoPJ0nE9PQcalW2s3KiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oUwfNAw+bWg5OBNk8/q6/no
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAnMZs04C9HXUfAVuhha+pcXmXi0cBBNzIp1U7i75hqCD2Iyoj+1tK/j2I16XSbL6C
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KA8irBFiq5/W4AZPCCvyETtXmXi0cBBNzIp1U7i75hqCBPvbRKR8thvzVk1X26jsuL
pZRe4QmM6mwnB4taJC3gHjgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAm4B3Ag2D3p4w7bSNc2ntyHmXi0cBBNzIp1U7i75hqCBXNeC+55xFSTR9M5uvUqnp
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAl3rLg6o85yqXYD++AAzpQHmXi0cBBNzIp1U7i75hqCBGaj768k10SN+yP5fo9B6/
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAh7hVnOz5PUBHuu2BlW1+f3mXi0cBBNzIp1U7i75hqCC//Rvc2G4pvSB0qJ5nWE48
JMu/mIob71FrLh75/bwN8jgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KApMLY1PcjjfSJ9uXb05pe5HmXi0cBBNzIp1U7i75hqCB2+MH/jZMfBZGAp2ilMks0
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAycyLZmANr31FpDWc84nQHHmXi0cBBNzIp1U7i75hqCDoJIeVS+iXRoEmk6vU/pba
1zV7SJMYIHpXwQ44MP2OgjgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAJ4xe4QlHxrcOE02p/Bz4vnmXi0cBBNzIp1U7i75hqCBbsF071G5Go/4IT9x8FLoQ
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAb2PYyGMm9wL+BfnRiHJFZnmXi0cBBNzIp1U7i75hqCDr0gOQCgqmRPWj3IAwz8Dt
2VE8eLlr40btFUWTGhzJdDgtCZJIAB9gvyW3A8wto8GDcJUeg7nTVihs38TkI9KAmaocPx8tshJHoaPL/9T313mXi0cBBNzIp1U7i75hqCAStGHJLv5uhh+RveuPMhSE
FJqAD3lIDMFTIw5+HZUauXiAhRj0OP4/9aXxYxMnqjTKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oUEtVciyPqWQFSM3qi1Jeqy
2VE8eLlr40btFUWTGhzJdI4R8zJhe3kc+ZAXe6nIBLZfV31d+TtvbkT3xj9q3UZFT0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCChfjy+OMgKKkHkisI7ivyC
FJqAD3lIDMFTIw5+HZUauS6ZpAk6HNlBMqLaF76l2TJUxpQyd0HAX6TAySxe+F5GT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oWOkBQiZxVTnH2HskJtjPgt
FJqAD3lIDMFTIw5+HZUaucpXYrIXimmZHNP1H+viUFjKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oVxneiYm0c+qWzgVmZPFGD8
FJqAD3lIDMFTIw5+HZUaufO8YitSLCzBPrjVtMeXNp8yzpinzexsSKNI9UWW2xEwT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oWtwoD+7URulgZOiPXUo1Nq
FJqAD3lIDMFTIw5+HZUauT4ahDUpcYnQwxk5FhqIX4nKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oWWsnG1LA+zQnfEQyZ4NP6I
FJqAD3lIDMFTIw5+HZUauWUeuGkpNoKLl3d9aqa9CpluPcqjj4KMfzKD264bGZmdT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oWqtR4gauQly8cW8igjMfXT
FJqAD3lIDMFTIw5+HZUauajgLvtWZIberlIDx4DJpllUxpQyd0HAX6TAySxe+F5GT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oU2HwmHqzVPY7XRyjNT4pJU
FJqAD3lIDMFTIw5+HZUauSclyTpXl4Quj6Q3Gr+y8/nKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oWQgjM9JmWijUB+uPFV78h3
FJqAD3lIDMFTIw5+HZUauUc0cHAHB4SzekJX9eHltf1UxpQyd0HAX6TAySxe+F5GT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oXL0dTF2jKu9PMrR9v7I8/9
FJqAD3lIDMFTIw5+HZUauVctGva8/AQY/n9QeqBBPbDKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oX7niyyk2qwy39hHnI9VqOy
FJqAD3lIDMFTIw5+HZUaucGcGijNHrIBqTN5nqcgxLluPcqjj4KMfzKD264bGZmdT0AdSo0+Ioxd3pOapgecMYKAnjCzmRrs+VQmwLFwhlVuFPQmZfjiIUgyskm+HWTk
FJqAD3lIDMFTIw5+HZUaudX9IwytLz07rTPwpptDmUzKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMYKAnjCzmRrs+VQmwLFwhlU9kAiChGUz9xvCdDzNSeYo
FJqAD3lIDMFTIw5+HZUaua4VLms5Cxlp7AMLXw10D3hUxpQyd0HAX6TAySxe+F5GT0AdSo0+Ioxd3pOapgecMQby2vpc1iIU3eKsbG/msDUGgyIc/DkbJJinnUgBuzjB
OChwhrvOT1+LtITHLffs5YiTzaeBQzdz2bF8pd5cNDLKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMRKxAH3sNjMnNXoJcwF2Iu4wzRQ/IEAu6lPvglUzIp4s
aJEFPP1T4G9Ta3LUsfD7iNIjhPUODMVs/IQDPrkR3NXKiCbRJr2HgYyrX3ljAm2I0bs3uyhPJXfV4SVgiJm4yHho0ig6M4VSzVM3SbAZ1acuRxZ4RKXNG56+mtoIEZxP
mCh/zm9/IK+Mi+eAf1KyA5LYlr3JANdr0phfV6F0O+1LF4omHtpUmYp6ePFaiTsts0LuJFF7bZuq6gp0PkAsIleS95MpjGHWW8qBzWZVpiPKiCbRJr2HgYyrX3ljAm2I
RU7c4+AcsoCp8kKEqxqyMgnmJKjU+EhcIjK4wmQbWitUBCseFF0+EF96SmKrurdy5lQ9WJAFsPmXNsjCcVLk3MqIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17
VIIOsWlTqOgtnYWIs2E9/DpBe9/O7ACRaRwSa4pynBfkaDyNsuEcIZXDMTTCnEuY0FDmPcE3UgPAVmunpzf9Y8qIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
DPaJ7Knr5nl/WXcA0ON4p1ablOdh7CRwTzFd0cpmXPhl8t7KD2TEUtwbRotsXcZQC3cSMVYQ5cb8vAJWDpOTQ8qIJtEmvYeBjKtfeWMCbYgSRqiVp9bf6hq6IpjBQBhW
7Wa14iv9WjgpVxqlnb2O0/Nz70gcCbxrQXmf1cJEJUlw78kcqjemwO5OHbioWdZs3tg36JZIjTN8D7VQ9R/VsnIHLql8/FShcQ41SVHzY3ZE9JWWoFQqmLP9vcmgPiAg
aWaRKigwaTE0ICP3dYGaW5E9DU1NvDtStEZIyxnvvAatCz9Gj6AYM4CjvJa1H0PYVMaUMndBwF+kwMksXvheRoEayJwYGQ9fRzfY+QWc56OCvAzcePFfFmnIty0uIJtl
UlGyf1c9ve6cNgns/mkd9rsDj0NuXkgIN52Huk9kFkG5yrCKAK4I/QRx7+aRjNkwMs6Yp83sbEijSPVFltsRMB58cROfMe6s7K9t/3ng+coK3f4K/SmYKkAjPch/T8NW
tc/k4BO9qK/2maGRQ6Nd1Ewa5kxf67wTtES6rinjigIyvZdw8hrgXJi4XeJ8oSnH0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNVDdEBUH1fBr0YhhKlapneS
IXF7fuEIbUn2+X510EUZmHJNA0U08lyz/1u6sDzpgbALD6FbEiXiyvwbK76KWtE56cdV+3ONhDnp7Kb9AzvcQokKJIyo56WBNXsbqnmq+U1Jld1HA3ixoQP+zzXD+t1M
gjL61U8H5kSH+Oyq/GhmLIJ/CWlu6LKGdJrNcWxkiatUxpQyd0HAX6TAySxe+F5GFdJkT329i7COnhM1KYxKoac5NNME6RdbdIjLB1avisew3w6DdcltZ0PdQN03ctb1
t8OKtKhX4CsnvTtgwKbQx2Sn9dj8yXDYuRCxZEqyw6lPQB1KjT4ijF3ek5qmB5wxPBMoSA+R/4beemn/L1nqhTeud70tX4Yhiuw78mHY8UvrZUD1tti+UlFo3ZVlGOlZ
i4LWhq7l5NwKcKW9iVpVUsqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFGGLgaDLcOU1AlDiD+2+8l1nRvHBbFnFTH8tyqXTcFkggzXQIqbuirq/jukl8QfiEN
8WP44/Hhv04wlArgTYQEocqIJtEmvYeBjKtfeWMCbYiqXU0HtT+eMVTl9oJBjZfXbIJTfYzg18hXY3JxSsFh4/UPbUsIXAkF/GvhyjcGTmWxugE/8w69wA1KCBKW0gCs
iZ+ne9XiMhN/TVmp7LhoAt4ER6ENG7m0FDD1bgBFTDorT0IBoL4Z0+hOhwgDG/l4GvyVY7ZpxbtZGnNJzEQiaJ0i7i/oG2GyKGGFH9fEMxXBVJ2dnbYdXE94x8sG5s+j
vdDEE33/Y/o79/QXczL/afXgIbG2KXL7lT6fOiJjyKr1t4TqmF+DK87kmRSb1CnqWZ+FADYvzl41DKotiIMvHevczVIjr21A+28dXJofnNbUfIDh8JQXVlNngfDy3BtC
yogm0Sa9h4GMq195YwJtiKuRCXjuaWzW1xmYO4DehHzjkzSQ6lswEgJAZleneJNy4pLvhU6uzGSsokiGnZulhQ3FwmP6lnDY1Y5TG118hrTy8WqfpQCtV86l/rdaJG3O
UxoQeWydCxDIplUUgtQSr/DuFpFTYUg8RVN19ERnN4vUJy66FSKqpKkQn5j2fqnSnb53OgZgTAwNdAbQ9KxKA9DyVbJ2SuORdP3O1ttCnIJqrV99K6Buhhy2PC9BzyTT
DT7g//IHiG2gW6jEeHDJCmT+OFExktJUgauPjekL8fDKiCbRJr2HgYyrX3ljAm2Iy5Wds1n057XZZv0gDvtT+X21ZbGXjVHjYYZGuG2ciqLmK9rf3LC0Whe+/aq12r74
cjveAzO+/7U58YwS7JUaF6pdTQe1P54xVOX2gkGNl9dr03PWdkO007tHX7mhMB2N+6yAqcur60LhaYAhg0929YTIWzPbNGKz92hyIJqibP0NgFGxPhBTHomBJZH6ns2I
5NjecheY3JPsioHKK53E61PVdLCKka7eyWNpSogHWBQpzJ/j8UjRrMeEErgdYTf4AB6QogYurEMhhBtyhsCrRlFCUL+72Mq/xOkhb4kCF8iO4kO5wWiofog8dGml4B4A
p650Ou2C1kIlhc1wkT221jNizoX/yZqyX0JK3BDZhs7UTS13V+Cv9nmqdg6nhaINlFJlcZ1d6MZaYjKKO/fbfalIzEz0vSdblY2KwNKp6M/afCmsSMQn8ESST2WieBIp
yogm0Sa9h4GMq195YwJtiPFevvcbJ018pnEiwmKnlurQOw4p87+FJMJxFDoeQu86y2ZmOBeLb2dpY5kGZGzj7vusgKnLq+tC4WmAIYNPdvWlV3fN3TgpaS0PsXSEL5HG
1qRdB0wNEM59n6HlciPS0MqIJtEmvYeBjKtfeWMCbYh3ezN5vKFyv1oKxzs51AAAyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
oFN7gHeT+ZseMhR+qjrtIqpr7fvUSRtvQlYo5wo+aeoc+TaNxDDi/A0Bd7t7rbQA5CJxF58DwuP+KzXN5XTAw+OstD6fvy60Dm0wiXjIwwBFtia/4eT5WLkpwWwiXSzo
l/f0pxG0tL91ifOD9P338FZpCiLBHtCAOfOolk5i0CXXXBAC6Vx2VUf6VLxt9KnJKY4HfTLQimKFPUOQjxlMMcqIJtEmvYeBjKtfeWMCbYiInuofpeo/KHrFqXBe2YOu
wFxnlphvA1QOZunS9R83kMCIGcCyY8y8RWVfZO39YK948byhxiKU0DE2C0fvggAyxrWiYC43u26AAWvP4zXni1ZWPo4SyGKZyoaK23bXbgrKiCbRJr2HgYyrX3ljAm2I
r7Cjglb1S1wPIp2b6oRPx8qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiIEayJwYGQ9fRzfY+QWc56OHVP6o0klEwO2A613MTJ8K
yogm0Sa9h4GMq195YwJtiG2aGZtJAW7/hBnchCAxhDj4bOSSMQ2D0BjrXvKwHbwmOvl+g4CKcd2n20BRSs17u8QyPFhrNC5LgmfFzqZ7mzRyBy6pfPxUoXEONUlR82N2
t+5ejgnMq6cFCUbL9uYwcQnAb4QkreZc8z0CyBkNBKZJld1HA3ixoQP+zzXD+t1MFQgud5e0U76HRqctBOPJw8qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiM0IMHlIf7x/msBKJ2C747PAiT5mGAj5ql4HQZUZ+5GA0iOE9Q4MxWz8hAM+uRHc1fdr2CFWnHLTtwVV42ElQ7NE2UmCDrBd4ywDS0YS5hqh
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYh9fAjVRLoLzOw+CHxUvqKrxr1lRClDItJoVOl4YU0eIWfgM2LCkO6jYV7LirKpNv8fRJxeMW51UrdpSJfv/5VU
gElHeJ4cHhlvjakLSzba1ZgAS//CDF9OepWJUNzoGTVNf3RUCPmzaE3QNwrVymL0uWYlo8vEGgrUtfVigxdV1DooEVAxespFc0Fkl9ViJzHd93Jg0pPUijZXofrfCAqh
yogm0Sa9h4GMq195YwJtiHRDKVZNP4lSwf13PICjvgO2YGUIPAj3YUTGRUOUqTTSyogm0Sa9h4GMq195YwJtiE2GJU8qPSq+3pj1a6aGi8oC6hxlxGIQn2yBxu8tXdq2
wu10agnpq9ybSsPW9UOYxTLhxmhYqgtFWuNBznYYsksefHETnzHurOyvbf954PnKU5Krw3DOjQrCP09JcW14dsqIJtEmvYeBjKtfeWMCbYj6la6pXbRlpgqIjQttKQ/W
7duPL00CTBnU7lE/7hcVRkCN/ND3XZvaB8pjXVLWrgPKiCbRJr2HgYyrX3ljAm2Ibcx9A3euJafUPZh7l1vZhcu6bpf0koypEhaaTKQKyZwz6tlPRqMfPuyLFxCoZQcD
eNHW4grv3qDmoS3a/SyIHE97jmH/NZ3VWrcypbH8BXk9byeZFLWBz5MiOduS6koFyogm0Sa9h4GMq195YwJtiEVO3OPgHLKAqfJChKsasjL31lT0h3gqRiP6OdFLVZyp
JgDFLYGPDrRF80Y6KUIGXSs4kPIiLKY8MdgYPltedM4bfihAz7uVEbgyCGk4GuBcVE8UNg3NkkHs5eb0lm1z9t4ER6ENG7m0FDD1bgBFTDrcD8dBQBgcZjBz164qcx/8
rLsCJ4obZeGMOmnz+7aU16zTfgvxC+rMcE8CGpf5qJOj9mc5nrVI/49F6ASK1RRXFXYR6m2Z6aZ0ZwD+pL++3Nski7v43HRpVdMY2TiLdzJmZicJwXgx5pHXyyvFB6lc
eZeLRwEE3MinVTuLvmGoILYMzw/JelQOwKYe0PdIp+PqtJB2Zua7duN3y50QepCyo94g30QmrHGoGHYKyrlhsoxLBfQTrASXbWueBcmb4PAWzehi8upxbgAPaVhV8n/e
0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+jRS6GUDc8782Nxr9qGJbkVsnsPmCil/eW3OJO5ycHjCuJIpgUq15Vb+ttxFlfaEQjT/QlWbTbsaIHkcd/f7edx
ATpTGK+P+Q1ZYdZpEjBom3IHLql8/FShcQ41SVHzY3ZE9JWWoFQqmLP9vcmgPiAg/qUOQozTq7BIjSo9+H7/jIiTzaeBQzdz2bF8pd5cNDKsOuI9G0DeFbW6PNFc1rta
SB6jnxB7C06R0m4uR2cisnWz2q/Aur74jf4b5HevAW6DcRdOfnzDCIY08vsxLu17VILgi9ptr6Yydmys3pc8wPGrnng6Zun0R29Zp9mK2L+m6W4Ih02GFZLFSFqUj73f
ittRvGrXOwvDNAqnrwf5Ke8TbH0p2sD6dONfI3aiD1htmr7Y5OuAcaxSnrrJ2SMT9eAhsbYpcvuVPp86ImPIqpaxv7kDoH/JAIeYKIjSGqDRWKSqc5EX+h0bd7wNrMhn
nixfgtigoCDhUqrWJMETmnN3ZswiTnL5vuEAVUNfGNphUH4cYnVi5BLqCdqytzkBSJhpOFU3JEBDrxHqs9QEr6GOGRbTFlHiOvUQpjJMgs3boghLczu6210BaMiqe2Ll
XIA6IN7aK96lFqPI7XaeZmGZ4d+DExHMCHWqrQC/Mplot5FrUyUcA3N0Ufv2sU3Ll0mjURa8u6sIGUa7IOUHDcqIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0i
O/Yj+KGk8Net4czuOrnLG1SdgNgb30eMafXQXIQNIFxhZCVudZalMVhV9NIEM38aMbFH5DJLyjvJpl+mDfB14p4XOUGOeKAXzu3Qu+KN+CxU44XP7LbQ0qpM+SrH2CV4
fUgoSjZJ0mfLOvTfraoVzhoZ5pG2DAwVL0uITmd2OLbKG/YMDHqG0bavCISZaX5lDWud16I4GcHq3rhoNGlTOch31/dBLbvgv0cVkpmj0PLGdJfhvVBy9rSjrrYYxvLr
ZEkljiuTsidH93CjhXspEImvX5jRYBoyP+S0/fQvdRoCVcPk9kgrpkZpid5xvrmyYAyEzu4aubwXNbGVPKkCDFum9ZySdYSfXfyudTxUmWsFK04fBmDzH2IzsziJx60F
EGeCych9GdCzRBY2uZ4wdHFTQ0gcvXqvk1d7T2wkurdAyaqwkAgzq4ApJkwTRqQMHoi6QCNavt+GRKi0P79ukKTHZL4OGnj2emdHss8NHCLKh/NRr0H+MQbvzML6s6p0
sNzzuRNBnsXJuVOgboO8msPQBkTlC+GCjDpyjgII7nJUhnv0Y0xKs+KegW9SjidpSeor+1VsbbG5l68CKHhk0kcuQWL8VUWKOqV9t0cIJdehpcyv7sO6Qv/zZP1yTR/A
txkHFeiwoR8H5V6zDA+GKjpFaV9ZjyW0vKCFXl3gH2+/8dVuvtoif0uXbkK8XoC+xlixEaAG3kWLAToVwmaNGxXSZE99vYuwjp4TNSmMSqFHX5TjNYmoUQ8w6SEjgQKm
yogm0Sa9h4GMq195YwJtiE2GJU8qPSq+3pj1a6aGi8oC6hxlxGIQn2yBxu8tXdq2HYiKI61yUxLtYKELLQcmmPusgKnLq+tC4WmAIYNPdvUefHETnzHurOyvbf954PnK
ijOWUChrMN/lu5grUNssn8qIJtEmvYeBjKtfeWMCbYjSJSRWN8ciwQ33PVyO2JPQyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
bcx9A3euJafUPZh7l1vZhbuMyCdiNemtp/TcvKy3nR/KiCbRJr2HgYyrX3ljAm2IyUSlwwO/0SYEzrRgH+b/2h7SS2uCwgZP0KSay+QnUSHeNRZSoynPMcnFCsa8rOqk
lmJwqSxzcxgAuF0utn7RHm4TwmiYB0JoXeD1l/zhSBmQOleJa9Vhtgi8KL9Od8yHyogm0Sa9h4GMq195YwJtiDW5eK8qFH8SxWA99ea9x9Fd383aHFG8pLoRz/CmKgF1
EJ0EIjq6xJOnd7qRumUKq5LFQhMGEKnU7caAyEG8+R0rT0IBoL4Z0+hOhwgDG/l4gx/aWa8EC31sKDj3aJX07cqIJtEmvYeBjKtfeWMCbYjqyOR6taVFkqz0FfANWuBp
CL0lFgs+zy6GkVajyRvIAiQPW4ye2H+zGKMNZOXtGj58jwzRHcqoavpwcxe2RLN5PBMoSA+R/4beemn/L1nqhZ78egxR0JnjSaLYxQyLSALKiCbRJr2HgYyrX3ljAm2I
GeY595iQRo89RRDbMJ1tCjSxPFJzcVv4lAwB0CeOj8nl86uJw5gW1jrjD4MYUNRdJx7JHwfULrDpdqo6GODMdpI3DT1waeDxQLTO5qtyfNWTFVjBEQM2FYQoCvNzCMLO
yogm0Sa9h4GMq195YwJtiOlCxOFOUT2VUhzEB8oO1CNtMaIY0s0bPLYSxF/sPqB/GRClyH9/Btolku34i8RSKHIHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+R
drPSVDp4R4N+iUp6b203PsqIJtEmvYeBjKtfeWMCbYiHOed2Q2nXBT39iI5kny6sIAfFXjDjb8IaS693+SRdxjzJ50rfYojBHGhbaKLEsPKDcRdOfnzDCIY08vsxLu17
YCTOfwZhQld+5mOO+u7zyNp8KaxIxCfwRJJPZaJ4EilJld1HA3ixoQP+zzXD+t1MM80io7RcGOSERyLZKJy3r4fPnUocYhLdJQeboMcSy2melWAGd8ZpgT5HRsec5BNx
NmWWg12F12lg4BpNV1U8x17FplJi9Rp+9i5hvBbZ0upw70Un1Q9IUc6G91GseXXAnixfgtigoCDhUqrWJMETmlz3doqaMwzLBtQ4hrh7jYfKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUaE9IrgBMrOk26YYKa/0V43lFTcqtgEDw/ZLyQeCYzrKWGZ4d+DExHMCHWqrQC/Mpn+0T2IRNcSxDgxcor2opWG
WVjmuB5r0rI62RBLMRyRXvNcU1RGB/yOhfm8ZosvZsXpx1X7c42EOenspv0DO9xCXQlM9Jqz3duOGVnCkFiOfaKrhBwMnRqV0s72OEmFtPdhZCVudZalMVhV9NIEM38a
MbFH5DJLyjvJpl+mDfB14sCd3b84K5sCXKusIxcsYqoDkGSLe8kPx8VxMZfCNN+SfUgoSjZJ0mfLOvTfraoVziniWtSiDodynwfQi8EmUU0uYpGIjaUi7tf3s84xauPr
DWud16I4GcHq3rhoNGlTOch31/dBLbvgv0cVkpmj0PILEltCxBmX0+vYC2xxr1LuQSZpSFO2o1eAup2K2DYwl4mvX5jRYBoyP+S0/fQvdRqX7Th2zvGM5MlOqBh8wG2u
TX90VAj5s2hN0DcK1cpi9CF9S8qJPc4urFGpjMIHEApbue5yF+q5KlkHq2ZwPrQNyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
rI8BKYpqUokaQpEv6JSn9cqIJtEmvYeBjKtfeWMCbYjKh/NRr0H+MQbvzML6s6p0sNzzuRNBnsXJuVOgboO8mko4o8jcEWrLxpxAI3DNFqcy4cZoWKoLRVrjQc52GLJL
ql1NB7U/njFU5faCQY2X16vjo7YYO3ShwTtw3Dsz5YgWMVak/JQci1J/FJS00RGj+kluENl35rF0a9MjLSrZzEOilBiWmNQv3Hs9dsPhWUTKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiHRDKVZNP4lSwf13PICjvgPx4U0oUl6i6YSNIlchnsCKyogm0Sa9h4GMq195YwJtiDE9REGn/7KqhKEhSd4rGl+LYGtvY/Vs1h2pytLRB97E
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKodYZQeRTkM0U/Iyd7Kwa0Mn8qIJtEmvYeBjKtfeWMCbYjR0o7Chg5TIi9E5naoHmfq
u0A7EV1bdj0SoV9IymjICIT0enC+em8umcqWs5uPjWTKiCbRJr2HgYyrX3ljAm2IEkaolafW3+oauiKYwUAYVg6xdiDJ5e1UmFkwW5xqSNbKiCbRJr2HgYyrX3ljAm2I
26us1gdlc3z0A9Mfk41iisJMBRG3r3K7H+sBRixxseLKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiEVO3OPgHLKAqfJChKsasjJhW5UPl3iNZSexloK3lSE7
yogm0Sa9h4GMq195YwJtiMlusTKEKUjFL1Tl9tYzFwA5bBHmYOQtmQPF0Dbqccjsyogm0Sa9h4GMq195YwJtiN4ER6ENG7m0FDD1bgBFTDrcD8dBQBgcZjBz164qcx/8
9r21GyGuDPGCD7eWQSjt+8qIJtEmvYeBjKtfeWMCbYgwai1uQltRFwwuxCJdykhtyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhPQB1KjT4ijF3ek5qmB5wx
/rQ9Ex/pa7QSWd+z3Us57wnAb4QkreZc8z0CyBkNBKbKiCbRJr2HgYyrX3ljAm2ILtQTCSOcbFir4MPu+NMuRsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
0yGRnPZE1s62DA8g752IHDkBOskn/alh5LtaIXu29FHP45sqZ4YalKRdnWUMnbqayogm0Sa9h4GMq195YwJtiHVND4742q96scThYqRhSVvKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiEIh/urAu31T7/2UbZfSq+MgPxzbi5ySN3VcZZ4fQJlk+oZHaffkJg0+n28A1ycdIclOYxqr8MDWCSrgReAzM/HBez1LjUzah+Vvp0QQHT6a
1n76s1dp7hfCS4MJRa2ddMkKh+D3K3YJSN8zpkS7pT78HlCE51bxhyMdtFmmYmpjTLPeuT/nwR+NqHjRr29dqotga29j9WzWHanK0tEH3sSBGsicGBkPX0c32PkFnOej
CaHOtUnJqSovpxwkgN5W+FyAOiDe2ivepRajyO12nmbkInEXnwPC4/4rNc3ldMDDjwCqN4OYZvEfVGkCqweDt6WRnKhK+FRF8UcAIoQlSvDKiCbRJr2HgYyrX3ljAm2I
ql1NB7U/njFU5faCQY2X13B7O6nB2ox94EkPd/bndklAjfzQ912b2gfKY11S1q4DcB0PT9BrXRqvz13urvxCHpTclEhZAeSBh0Y/zJsKWbs0NlttMI/Mk4dF6gZ+5Xkj
yogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YWxGUXId7FQvysB6pbmHQe/sDoEcCFGKWpDb8rs6v+sq3EeRs8ohL2If1uJ6WG8a18HzeD5fVv/bQxZq07acXvJ
iuHdGjE3t3MBqu6uWezOgic/kQdx3MjegaW3tiTKEDN5l4tHAQTcyKdVO4u+YaggD8Lt/ykt2+ata7FGEh1AbSYAxS2Bjw60RfNGOilCBl1IVSkI7KbAY9btSsWgi6RQ
GFtblCiiDJ+LjPDqtqNYrP5Y0IrBpttDMmPH6IkfPmjizk8ZLLY+mFHmOXZl4WWgr3BHxdEdPsnrYsA3HT2E8EtthOIIO3yJR+oDaBaCdDIuCJQdxY6Vm/1C3HU3Ixmo
G+zB0snn9mpFcDFIqM6JDlyLc39Bgz9Qs1LiWKpiuwoK8AiKI29mzCpW7jADuviwaeNS4YONXZsffwku6s+5LN7TLRmxdYRpn9b++ETtzI/ijJr3D21a9bgoc/xko+/y
JN/taMPTlwBb1mlRZXmNmND+w5Q1xOQZr8clYQPdt3ExX1S05TxHKSYC2r8nd6hQ3QSvOqLoFAXr1LdrwTUjysNDtnGNeCDVoMISkOauPUB5Bou9cYQ4f1cyiuBfWpYe
RHl8A6pExkjxxo3VttEVlWgOaAhQA9iKo8bjTaScZBRImzE0t7W06yA/+OvXsfALkEhE+JscsAzzIEdqIdzL7hr/+uzQNRirOAhZ4rT2DmhU6co60/5xo+OxKJHfFKod
pDAixgPdhmk/Wm6tR3wtrPk7EI/U1i4rWutF5UXgsOyYGcXjFLDJBZdyRS85uFGBa4OqlpaoaCfs3nfliNoaS1GTyKMbnzxB6ULWAgKbZGh84z1aShWFrytHqdspJLuA
3A/HQUAYHGYwc9euKnMf/LGrzXUeizbA6eo+Jdve5G1WapOQ5OY7MWfmsHTheYcSS1VBvPirY4PczGpkxwLsZwsy5njU9VN9aUKRiXgVWnegb5NCX0h2/ImG4tzBlm2A
ENQ/ceEMamHXT39DPbMVmET0lZagVCqYs/29yaA+ICAqMUSjRvCzscdc7DAlYmnVyogm0Sa9h4GMq195YwJtiJGwSiYIsMKnaDIr3yqbIQimkBGFRbLCzLZIxQpeMr2l
yogm0Sa9h4GMq195YwJtiKGOGRbTFlHiOvUQpjJMgs3+Ae71lURXxklgq1G3aKLI1A6Y4zXqsfGOQk9PLoLFvdahIyIuQnw+ZKKHkf3lYD4EOHAYSUZrnzoCECeKvZtG
m9yqLWEv6hg7ZeyvGmM/erFSkEQchg0CCKwa0FlvnOopsBaa+693yKVXWJwNX13Lnq0WEosBAWqSs3pGqAUjm1SdgNgb30eMafXQXIQNIFxBHZ58I7/MXFr/Gna5HWtw
rzqys6hXw1zuIEwzpvo96DCPESMbaD+NVaJYQWhGtCTKiCbRJr2HgYyrX3ljAm2IFdJkT329i7COnhM1KYxKoTYHXYgL+ycDuhVAjc2Hz249byeZFLWBz5MiOduS6koF
XKdeucuWucS48SrzY1v4A90ERJysncLlt5pAkNIJoOxkSSWOK5OyJ0f3cKOFeykQyogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBntLhF5lk8tVI+Enocprf5J
N6XC52fW5cz7b62pCMp2A5DZ503Uvxih7GO+IiY0HXoz7KvbprV8XOBY069ySxyfYAyEzu4aubwXNbGVPKkCDNMhkZz2RNbOtgwPIO+diBz9DcI1aD0KXLqpOSiSINdY
ZizVc2/sA3Fp2ONaG7TyaQqOyhoKxJaGCt4myMNaNZK5TX8WR+PzrbowU/ZBiy1Dww5AaTDDLgt2hMsUC/7iQIIB70UJXDnhmG5lPX6Zw+M2ZZaDXYXXaWDgGk1XVTzH
wXs9S41M2oflb6dEEB0+mqqZqlinSfcSiJ+KmLr8CWxfzNlE3Ikc84dw1qUxGpu4MKDACeSl9X6kjJe6jBqOBJWPDLHiuTuEEDeIHI/VmgICD+Ub2TcuiMyZVl6wfe9+
fUgoSjZJ0mfLOvTfraoVzlfbz7inj2VIuy+kIhIle82LYGtvY/Vs1h2pytLRB97E5CJxF58DwuP+KzXN5XTAw9lCV0UafUhRzM4chONDFDDXB8Uw8kWzJK0n3Or9b9DF
yogm0Sa9h4GMq195YwJtiKpdTQe1P54xVOX2gkGNl9czMNcJlT5WkLsW1MKAXmaO2IxgPx4X0/eBdEw8eySRiND9c+27Zzqo9DEnA6UkxcqYBV5I8BkV+lB2oSVXsQFg
zokdfAWKlXjJHMWLsHayocqIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mF7+YEhuq6iWrme09aV3SWG8qIJtEmvYeBjKtfeWMCbYgxrbnphwwLSgvsTZlRprWB
Cez9tkRYYayMYcShU4dsgi5ikYiNpSLu1/ezzjFq4+tPQB1KjT4ijF3ek5qmB5wxPBMoSA+R/4beemn/L1nqhTa5zmDY57Uf/npYSekQ2dlE6ICSlzr49ovY7MAV/IEd
bNXYjYq+HulXNX3jjw7U04xLBfQTrASXbWueBcmb4PCXfuDIEmEwlORSfimFsDnfg3EXTn58wwiGNPL7MS7te43SQmvmCzEG7Ealf+1WqB3+WNCKwabbQzJjx+iJHz5o
qQQOfH6c5lWt2+6sW62jCKoTeKc3MfpwxlYlT8b2xwzvE2x9KdrA+nTjXyN2og9YX34wyo1hWds9VDBa1X6+CunHVftzjYQ56eym/QM73ELoCUJ/yXPCpBCp3Xouux3f
CvAIiiNvZswqVu4wA7r4sI7iQ7nBaKh+iDx0aaXgHgBbzQIbnjnQSeLTnCw1O2W/iqufVS6TOUhCNpjOJbgnTt9AyWEX2b/RNsThBZZLs/VAyaqwkAgzq4ApJkwTRqQM
VBFsixLYh2WHxWyhSqoQQ8A4ozyAV26NeSuwgZY8b2DikrYJK2etvaGW8ZwfCAr/tpSNOhVcLO0f3tJptFHxFipyDAfSnH2R1flpgIjDhkFhf4iAA8hLomP+1mbfh/Ly
HnxxE58x7qzsr23/eeD5ypjQ0tiuNAp9szp9dU/l8SXk0VS+9C3ZAyXzn1yGFd6Lx2aYVm8+gMihdStS3dohvwFWJ4YrzczUJzWRf+tmTYOEb6QVL5xgZ91wIrUIn2GG
y4vb+EDQ8arvuwunp+dcYytPQgGgvhnT6E6HCAMb+XjvE2x9KdrA+nTjXyN2og9Ycjrg2djo1TimXlYnaDFobJ+Kj9zJBmHwnwr4b+bNQXoVdhHqbZnppnRnAP6kv77c
k+xUP+j7FAHOojBCerLIHHIHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+RoG+TQl9IdvyJhuLcwZZtgOXN2D8F0byLJ4Akjo1vFWORsEomCLDCp2gyK98qmyEI
SB6jnxB7C06R0m4uR2cisgIP5RvZNy6IzJlWXrB9736hjhkW0xZR4jr1EKYyTILN6Whyzlz2OamAnp3FuJ1xcdp8KaxIxCfwRJJPZaJ4Einw7haRU2FIPEVTdfREZzeL
yt0OY2aNKH0mhkBxBvC15J0jLuJ453UF9sDIOBJ4ZJPKiCbRJr2HgYyrX3ljAm2IKbAWmvuvd8ilV1icDV9dy0mEg2D7stHPgYRi2x3I6w+xUpBEHIYNAgisGtBZb5zq
QR2efCO/zFxa/xp2uR1rcNcADDE1d7OBQbq3lI0FoDkCeZlAhPUv6FgP1FwivFOXyogm0Sa9h4GMq195YwJtiBXSZE99vYuwjp4TNSmMSqEQV+3xIzO0JwUMQ9jHkIce
yogm0Sa9h4GMq195YwJtiFynXrnLlrnEuPEq82Nb+AOLWFW1UKCnZIIhsdfXRXpLTkKvadyYY9/dnJDcHdolicqIJtEmvYeBjKtfeWMCbYhFTtzj4ByygKnyQoSrGrIy
/F7fKz9nsDQCTNzTNI5AP3JjQqQZ41m7EFvfmrlGJQGyXixi48mGtaG2s5ovbtuU6QT7C3PmFwdTYe+6LoJGCTpvG7Rq1BIm++JChRdCpTPTIZGc9kTWzrYMDyDvnYgc
uc/k+OXiweAW5ELnA4Vm4Loyquy2+YsYeXBvirbGNgs9bO7VZXP3hxhO7ddihD4V7IfcRxofuyCu3Yx+7uFqpPFEnhS83uXIE5iwxjRbKTKn3pbdW2cgLd+9aiKk7ztC
9eAhsbYpcvuVPp86ImPIqoAfarH8HkvbJa9S3vH8llp87WfP8NVMT6t68FK1JcQ7Ko9m9Kwl+fV9EHP8S9v7iiW6zJk0so/Z/kO8I07XoVqfHGHWXpSTo7z0ZoJIsD00
Gv/67NA1GKs4CFnitPYOaIEayJwYGQ9fRzfY+QWc56NIdtkISh2KfbL0NSvgQdYXBoytnJAlkhAUaJHvWi/jRuQicRefA8Lj/is1zeV0wMO9hX3tY7DdCBs0O0A8+JXS
tgS7lVXpG9F8pfSLbLf2u22avtjk64BxrFKeusnZIxOvVz6gH62yW0/Tj9EXkQKUcYiq+rhUYKHxXdsrJjOelXjQTgCEN7leBE4lrpouiKFxruNlKVzC2NYn40hNrnNQ
RSlGxml3XWzK/L4AwcIEJU1/dFQI+bNoTdA3CtXKYvSYGcXjFLDJBZdyRS85uFGBa4OqlpaoaCfs3nfliNoaS8g3sMrtZZ1zMOlf3tLV4p3KiCbRJr2HgYyrX3ljAm2I
bcx9A3euJafUPZh7l1vZhdUGrVW5YS6Dd3/yXK9l4wnKiCbRJr2HgYyrX3ljAm2IeNHW4grv3qDmoS3a/SyIHB8wa46o3Eq1t+ONB0ds4J9yO94DM77/tTnxjBLslRoX
yogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBkj24CgSt7Ek3M46qp+eBRwyogm0Sa9h4GMq195YwJtiLziLrYXES/CFG1ZCH1SN2U8iMs7LHNqtdzVo0Jm9XJT
JBfXb6CNpgIE1HlBywlXSN4ER6ENG7m0FDD1bgBFTDrcD8dBQBgcZjBz164qcx/8savNdR6LNsDp6j4l297kbTPq2U9Gox8+7IsXEKhlBwNLVUG8+Ktjg9zMamTHAuxn
yJfLoc89PHHBPt6rH1j7f2e0KmmL/S48dP2BLR9cPkX7ZondZc3zWM+wDjA41I6CeZeLRwEE3MinVTuLvmGoIA/C7f8pLdvmrWuxRhIdQG0mAMUtgY8OtEXzRjopQgZd
SFUpCOymwGPW7UrFoIukUD4yY54mHwRizXYph4BUepT+WNCKwabbQzJjx+iJHz5ouvYviyBRLiSbYIKbsftQzvNLNbtjqh2E5tBXf9jKf+iYD/WdU0fQEptj8s8V7By0
rNN+C/EL6sxwTwIal/mok+eyjcHGEigc7zLy/sRJUImjbf4MF/0/CXFqlQRluXZWYtkSFpHWmUPN9F8o8AN7KqPvFAbwZmpsLpIQca621GRE9JWWoFQqmLP9vcmgPiAg
IAKDWCFOwDcDiXTtFLd0leq0kHZm5rt243fLnRB6kLJtr9X2t59oVCVgPD+TiRi3U0ycmPalEGnIcCRilCOqnipyDAfSnH2R1flpgIjDhkEHfc6gwaodS/rASaXSxs16
r3BHxdEdPsnrYsA3HT2E8NFLoZQNzzvzY3Gv2oYluRUQ/QFWUWPHS6zQYNWUye1nG+zB0snn9mpFcDFIqM6JDok/lomcbCg87NFE3kCDf0qoO47DyXYZ/rK/4lGYa3iG
RP5WgZpjjT10r/GxJyAbAcF7PUuNTNqH5W+nRBAdPpr+pQ5CjNOrsEiNKj34fv+Mo0bMpnimJzvP4DGDxhMlvvweUITnVvGHIx20WaZiamP5yszANBwVz+1JELSvmCeN
Il1Nvb57nXfyN60du1Io6DQkEy63pE+g3elHkjglavRC78hPCHOnebdjSN7gozVd8aueeDpm6fRHb1mn2YrYvwJFjksBYgk1p6QmOkhKC6YEOHAYSUZrnzoCECeKvZtG
xfks74RvMWMyhkptSVSbhMZYsRGgBt5FiwE6FcJmjRugU3uAd5P5mx4yFH6qOu0iD+OErqmEzktaX7yoVmkpmtFYpKpzkRf6HRt3vA2syGdhZCVudZalMVhV9NIEM38a
XCaHntcoy8MWPz16fh7i0ioxRKNG8LOxx1zsMCViadXKiCbRJr2HgYyrX3ljAm2IfUgoSjZJ0mfLOvTfraoVzohzv8UttRhCdquEfRg8zMxcgDog3tor3qUWo8jtdp5m
dtlVJX7Ir0QL1NYIDikGKpH5Z6TamolI6pILnW++Ez3ytPuUgchKkGh2NWQazlaN2IxgPx4X0/eBdEw8eySRiCmwFpr7r3fIpVdYnA1fXcuerRYSiwEBapKzekaoBSOb
VJ2A2BvfR4xp9dBchA0gXCF9S8qJPc4urFGpjMIHEAqvOrKzqFfDXO4gTDOm+j3oMI8RIxtoP41VolhBaEa0JMqIJtEmvYeBjKtfeWMCbYhAyaqwkAgzq4ApJkwTRqQM
sqX9wTkWfLIFmYB2lI8Eocob9gwMeobRtq8IhJlpfmWBq+4lTzGwwrsjFrZ/RxhvhOUyQ4iL1rrhSytemnzIkiHiIPGGXZ0wMXj8mh67v81Mv+FRuDwWS35pftzEc+0a
ql1NB7U/njFU5faCQY2X1+B51wQZFsbrRzV5rlNwAKRgDITO7hq5vBc1sZU8qQIMuWYlo8vEGgrUtfVigxdV1DHeQyUVwiYqY8nauQP2mnBqBR17tWQpht24Vd8GxHAh
3tg36JZIjTN8D7VQ9R/VshXSZE99vYuwjp4TNSmMSqE2B12IC/snA7oVQI3Nh89upMdkvg4aePZ6Z0eyzw0cIuJZtZ1ZTnnSclH6ET18z+zdBEScrJ3C5beaQJDSCaDs
th3t8qtYNrvSQOYPseS/smOLKN/NVM9esVtn30j64skefHETnzHurOyvbf954PnK3hsqQLJ275uGgYBZf9Ulk6GlzK/uw7pC//Nk/XJNH8D6la6pXbRlpgqIjQttKQ/W
BONagr2PcZ9zXBKBZWw6Od2cUX+kBd2DoV0AjK3UdL3KiCbRJr2HgYyrX3ljAm2IEkaolafW3+oauiKYwUAYVkZtPSwSXNl5c/iwZVNtE//KiCbRJr2HgYyrX3ljAm2I
eNHW4grv3qDmoS3a/SyIHJz0zE1BFXlYc9e+rEK4o/n7rICpy6vrQuFpgCGDT3b1yogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBknAU1R8znw7bPIEQmihd+3
yogm0Sa9h4GMq195YwJtiDW5eK8qFH8SxWA99ea9x9Fd383aHFG8pLoRz/CmKgF11pJ0rhnlxI2gt3W1jwhEJd4ER6ENG7m0FDD1bgBFTDrcD8dBQBgcZjBz164qcx/8
Ph0oOoLhEVQM6X0gGd3iKsqIJtEmvYeBjKtfeWMCbYij9mc5nrVI/49F6ASK1RRXprRwCOACWsY94xHlL088OcqIJtEmvYeBjKtfeWMCbYhPQB1KjT4ijF3ek5qmB5wx
PBMoSA+R/4beemn/L1nqhTa5zmDY57Uf/npYSekQ2dlE6ICSlzr49ovY7MAV/IEdo94g30QmrHGoGHYKyrlhsoxLBfQTrASXbWueBcmb4PCXfuDIEmEwlORSfimFsDnf
0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNVCDY6kpPPo85HB198p+T1VPWzu1WVz94cYTu3XYoQ+FeJIpgUq15Vb+ttxFlfaEQjT/QlWbTbsaIHkcd/f7edx
wvJPdEp4FyD7l8NphrAXxHIHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+RiqufVS6TOUhCNpjOJbgnTkHgeuOxDcblvjNo0qQTZVKsOuI9G0DeFbW6PNFc1rta
SB6jnxB7C06R0m4uR2cislAU4bEI5ktLq/lx1MzGeZODcRdOfnzDCIY08vsxLu17jdJCa+YLMQbsRqV/7VaoHZ/5JZYlSzIWeUYgMrSqKrQfiy7BRnETsWsNaqMWIHVT
ittRvGrXOwvDNAqnrwf5Ke8TbH0p2sD6dONfI3aiD1j9QHt/1z9lEtaQRKL2awxsNmWWg12F12lg4BpNV1U8xyv7Z5piUGdNYHFs6eY1Y73hsgeBRaLW5blz0nv6+dao
nixfgtigoCDhUqrWJMETmvqEzQZwm4zRhJz3DndtCS45OXkyxINhjaYTVCPopW9vpx6joFOeblw1gjdWHYnG7KGOGRbTFlHiOvUQpjJMgs1CsQW5q4MhKtZrSXHYjizn
sECBbdgdd4Jyfk9VZ2LW+GGZ4d+DExHMCHWqrQC/Mplot5FrUyUcA3N0Ufv2sU3LXys6JsSdYbZbRp0UbTVL+G2iUvgurAN1etzYyDnz18Ppx1X7c42EOenspv0DO9xC
6AlCf8lzwqQQqd16Lrsd392cUX+kBd2DoV0AjK3UdL1hZCVudZalMVhV9NIEM38aW80CG5450Eni05wsNTtlv6Bvk0JfSHb8iYbi3MGWbYDlzdg/BdG8iyeAJI6NbxVj
fUgoSjZJ0mfLOvTfraoVzi/I2KEtDlbR8rxBCDCPxoGLYGtvY/Vs1h2pytLRB97EDWud16I4GcHq3rhoNGlTOch31/dBLbvgv0cVkpmj0PLGdJfhvVBy9rSjrrYYxvLr
2nwprEjEJ/BEkk9longSKSmwFpr7r3fIpVdYnA1fXctJhINg+7LRz4GEYtsdyOsPsVKQRByGDQIIrBrQWW+c6iF9S8qJPc4urFGpjMIHEArXAAwxNXezgUG6t5SNBaA5
AnmZQIT1L+hYD9RcIrxTl8qIJtEmvYeBjKtfeWMCbYhAyaqwkAgzq4ApJkwTRqQMuyaF2Javi3kp2JjLlCaGyS5ikYiNpSLu1/ezzjFq4+vKh/NRr0H+MQbvzML6s6p0
sNzzuRNBnsXJuVOgboO8miPaUpFzumFWWSogY9WCAAtBJmlIU7ajV4C6nYrYNjCX0vZ/C5D4uxV8hGR06yAxc+pKep3K4KKr1fcrHssd1vxcNTOtCc+GcEoyWXd2sbju
txkHFeiwoR8H5V6zDA+GKjpFaV9ZjyW0vKCFXl3gH2+/8dVuvtoif0uXbkK8XoC+l7Cgg+em/nfKS7j2BBT3FnRDKVZNP4lSwf13PICjvgNt7grx43jnU1T+b+AKf9UV
NJcVnl8nC2lJnazY7jtP2U2GJU8qPSq+3pj1a6aGi8oC6hxlxGIQn2yBxu8tXdq2q3Ls4y1uxab4Yhmf9Y+H3afelt1bZyAt371qIqTvO0JU6co60/5xo+OxKJHfFKod
uelAITd27+eTX80priqeGuTRVL70LdkDJfOfXIYV3ovR0o7Chg5TIi9E5naoHmfqu0A7EV1bdj0SoV9IymjICPYlg31LNpf6Qho6eSE+V7gEWzcW8X/s/esqwkM0mpq/
bcx9A3euJafUPZh7l1vZhfDJkwYq8v37bjcG7XMu4JVWapOQ5OY7MWfmsHTheYcSyUSlwwO/0SYEzrRgH+b/2h7SS2uCwgZP0KSay+QnUSGN1lLHmEziY55ufOqahEJM
071Ryi+qiA0Hhdug1eNnNrrgGdsgh0doAUAlFSabW/HxfHSD+wSWupUBddgQ+1+5sf1mjBGjb/lplAUZ7gFi+ZLYlr3JANdr0phfV6F0O+1LF4omHtpUmYp6ePFaiTst
F5SHyKoQleKKaKVr0jBH8Dwzcn5SNp1050nFAtYxwZnKiCbRJr2HgYyrX3ljAm2IRU7c4+AcsoCp8kKEqxqyMgnmJKjU+EhcIjK4wmQbWitUBCseFF0+EF96SmKrurdy
In3CToqLskqBJ9JnitW/9ew5oHY7Y9hT51NhYA050NCDcRdOfnzDCIY08vsxLu17VIIOsWlTqOgtnYWIs2E9/DpBe9/O7ACRaRwSa4pynBfkaDyNsuEcIZXDMTTCnEuY
VIu5lQpfVlhwwH/MkzCs96VjCWUq1lGm2UiZV2CVqsUpsBaa+693yKVXWJwNX13LDPaJ7Knr5nl/WXcA0ON4p1ablOdh7CRwTzFd0cpmXPh6umXiJHqqRYVxh0LT6KtG
k9XEv/OF7LYZp+Mcot0JjMqIJtEmvYeBjKtfeWMCbYgSRqiVp9bf6hq6IpjBQBhW7Wa14iv9WjgpVxqlnb2O0/Nz70gcCbxrQXmf1cJEJUn6pgYt17pkmx8wU3mToX/F
eb9Y1CanRI4TrADaCSAu9XIHLql8/FShcQ41SVHzY3ZE9JWWoFQqmLP9vcmgPiAgaWaRKigwaTE0ICP3dYGaW5E9DU1NvDtStEZIyxnvvAYVTG2mWSIVB2yZMPpf2du5
SuRgEPcZNWUXRsTWxU3aGYEayJwYGQ9fRzfY+QWc56OCvAzcePFfFmnIty0uIJtlUlGyf1c9ve6cNgns/mkd9hz7ocyWY6xBBQ2jUWsKP7QpgowpcDQ4wwuGNgmbTUsU
yogm0Sa9h4GMq195YwJtiB58cROfMe6s7K9t/3ng+coK3f4K/SmYKkAjPch/T8NWqmlUgV25a/mU7ZlpoFzxbULXfb/spnUIgIXBGnLGTUKbGD/qhaoVsQxNXv/sH827
0yGRnPZE1s62DA8g752IHJI3DT1waeDxQLTO5qtyfNXeEqvtTUBiZb66oZmBpyNhsrh1QWjW5V0j+Ti0f12k3haATFz8Bj5Pq6sT7vfisEm2F8JTI8fckIfUO9H6EUKU
6cdV+3ONhDnp7Kb9AzvcQpw6hhU/Mmkfov7pQ/LGNtiyclL/rs+tsr2Vlo2+g0Qjhc4jSwzDsq2W8fvr8FGgKuYQf5qmth57HmMpVhfZb3vKiCbRJr2HgYyrX3ljAm2I
FdJkT329i7COnhM1KYxKofEY0+d/flzq8HQ6cUSkltsiapC7PpNOCu2aOu6tZDMpUUNw5O9HSCTA/bZqqQWJeJzc6TfRDiWl6NCjnP/VxG9PQB1KjT4ijF3ek5qmB5wx
PBMoSA+R/4beemn/L1nqhcdwOw2mT9ttauUpvtQ0jR7rZUD1tti+UlFo3ZVlGOlZrBnA+dBWU1MLwKn6BKiQaNiMYD8eF9P3gXRMPHskkYieQ8QsxJAEjcphVGeA8TFG
qJI7YEbeIAYkNBFAqjXCBFNJTmUAjnbSeteKmu9tItyudynD0odqE1YjrinIp7KOAYklrXzFCNtSC4n/fPf2VMqIJtEmvYeBjKtfeWMCbYiqXU0HtT+eMVTl9oJBjZfX
ayx+TXsHKVcIeVkxag3GCvUPbUsIXAkF/GvhyjcGTmXJ7OQw929ijH8IssWq7utlaLPYK/qqLL4WxNyYQ/Hnzd4ER6ENG7m0FDD1bgBFTDorT0IBoL4Z0+hOhwgDG/l4
+VZn+AKvy9ky1zD8ks0mxp0i7i/oG2GyKGGFH9fEMxVCm3iXnG0Is88Y7YqrIlNDSuRgEPcZNWUXRsTWxU3aGfXgIbG2KXL7lT6fOiJjyKotOAzdk3Fu0STcvCDdr17U
WkkXKG6MR8jekvo25zyGsuvczVIjr21A+28dXJofnNYi0I1PyTTwXDq7XBBqILbvyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60++XatWDphohNdferUtWvnGR
SxeKJh7aVJmKenjxWok7LXvGoJQ1WiUdvVpjSb+nj4twXT5xM79Jwh4xO8iQFjSIyogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBnJfO2LL8f3izAKiukYtaxS
3Dv/kXzwIqsHZNfuHsRwxgp7rJy22YbSdtKZ6GqRSXJmT1CGmPJ5xxBLbM+dnreXg3EXTn58wwiGNPL7MS7tewqYXg0Um8YrYAynhIuHLAiA3z1H8CtDPtBxz7TSxHvi
B7T/3l3ivpLfvRrqHqOJTOuyPncPwSUUFUkiRkCJHTzKiCbRJr2HgYyrX3ljAm2Iia9fmNFgGjI/5LT99C91Gu9/hiNFCWR9Tb6YBd57yWY85SqxfJOZ5yMgRDjKslEE
LnBPLbCjOLf5W48WzrdlRwRiEJWN3PTM0kll+sZ16//KiCbRJr2HgYyrX3ljAm2Ibcx9A3euJafUPZh7l1vZhdwwHeP9GNTudovgxYe5DsvVia9Tqd40SXXFLd6A1m7g
dgOsIkItmN+KKZz9CdIJfNzB98jR0TzjJrgFdyQttTNyBy6pfPxUoXEONUlR82N2BgFkoZbbTLQ27IEut7gPkVm+QyoExqG1bOm849l6BxxItcTvA2A6xlY4KqarfLp6
6w8xhrewvxm4YrmgVEpIM5ZicKksc3MYALhdLrZ+0R59SChKNknSZ8s69N+tqhXOn9jKC3NjT5Dohtn/6/uoVbBsB+/EoPvXoFhkTYyqxFsc+6HMlmOsQQUNo1FrCj+0
JPF7e+72CEp48EcdMPvgYMqIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKod19aH7cePAq6MZbC8SRQDENanX4XjZtFlnLC/eFWfMYutE6ixkwHSeBeuX/b+Jm6n
pu2Et7bm7cQbNLRq0Vl6u9MhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbgXVHlH7eFefep4oUREe9g3bK4dUFo1uVdI/k4tH9dpN6x1k/geE+a5KXIDjt9vhnu
thfCUyPH3JCH1DvR+hFClOnHVftzjYQ56eym/QM73EI2ync/VeD5h/PmN1qrYUcTsnJS/67PrbK9lZaNvoNEI4XOI0sMw7KtlvH76/BRoCovQEwvdSQHgqmlpT5UkMlb
yogm0Sa9h4GMq195YwJtiBXSZE99vYuwjp4TNSmMSqFrrpqRkQ+d2h9d4h4bOA8GImqQuz6TTgrtmjrurWQzKXhsveimba+8ycR4KJvfvjmc3Ok30Q4lpejQo5z/1cRv
T0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oV/eRn1DsV5jcaRK9CvTvbM62VA9bbYvlJRaN2VZRjpWYsuNQlaNH9qRfRR/sbFDEnYjGA/HhfT94F0TDx7JJGI
nkPELMSQBI3KYVRngPExRkqKnJqxJ2neuVBB54fzCERTSU5lAI520nrXiprvbSLcrncpw9KHahNWI64pyKeyjqJ1CU2I6staP6HqsSDhGBDKiCbRJr2HgYyrX3ljAm2I
ql1NB7U/njFU5faCQY2X135mhxZX9yeEkbTvCkuSjlL1D21LCFwJBfxr4co3Bk5lhoZlICPJIv6ZsTXmOWnFgGiz2Cv6qiy+FsTcmEPx583eBEehDRu5tBQw9W4ARUw6
K09CAaC+GdPoTocIAxv5eEevxFXqJ3noznTLpycdOS2dIu4v6BthsihhhR/XxDMVeN4YgOAst2EimMJ5oG337UrkYBD3GTVlF0bE1sVN2hn14CGxtily+5U+nzoiY8iq
exITj1J47G5Svhapp2Rg5lpJFyhujEfI3pL6Nuc8hrLr3M1SI69tQPtvHVyaH5zW+8f3BVp5B+Lcs/Zn3xwmCMqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
cu7alnr7V2aeQr2Yz96HNUsXiiYe2lSZinp48VqJOy17xqCUNVolHb1aY0m/p4+LPiPXOajsbMeVJOJ4tRrVOcqIJtEmvYeBjKtfeWMCbYhuE8JomAdCaF3g9Zf84UgZ
iRo+cZqFjlF6K2nSqKrhTtw7/5F88CKrB2TX7h7EcMYT0a54sENZw+jybA7dRJyqZk9QhpjyeccQS2zPnZ63l4NxF05+fMMIhjTy+zEu7XsKkGCXziHgzEngnMzTk8Nu
gN89R/ArQz7Qcc+00sR74ge0/95d4r6S370a6h6jiUwDCfLDeUYFvtgw6pGmaRcxyogm0Sa9h4GMq195YwJtiImvX5jRYBoyP+S0/fQvdRqaZg1WlDnPQpWwHqClaaYz
POUqsXyTmecjIEQ4yrJRBC5wTy2wozi3+VuPFs63ZUekYohxx+3U1Fu2dc1K+jcTyogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YUF/lsays5qbnPAt2s3ThE+
1YmvU6neNEl1xS3egNZu4CdeETDc28GkSGEZwHlniG7cwffI0dE84ya4BXckLbUzcgcuqXz8VKFxDjVJUfNjdgYBZKGW20y0NuyBLre4D5E/TEJN6HB83a7O7YVmDK2z
SLXE7wNgOsZWOCqmq3y6epTI2S6t7SvyKjVoHnuVyZGWYnCpLHNzGAC4XS62ftEefUgoSjZJ0mfLOvTfraoVzmuBZMhdVo2J8OCMsNLkqMewbAfvxKD716BYZE2MqsRb
HPuhzJZjrEEFDaNRawo/tDrb6aU159MSDqURtJgR0uvKiCbRJr2HgYyrX3ljAm2IVOnKOtP+caPjsSiR3xSqHXUTaGrmWxoH+fP/h/J4XxLWp1+F42bRZZywv3hVnzGL
QLzQXU7AJsorsdvoIIPwlKbthLe25u3EGzS0atFZervTIZGc9kTWzrYMDyDvnYgcuc/k+OXiweAW5ELnA4Vm4EZBBoH27j54BAyNGZCM/d2yuHVBaNblXSP5OLR/XaTe
E0l076BJBMSNYVceFQKKPrYXwlMjx9yQh9Q70foRQpTpx1X7c42EOenspv0DO9xCPDgUBf2JruebuuiRDh8RkbJyUv+uz62yvZWWjb6DRCOFziNLDMOyrZbx++vwUaAq
Y6JdB5GQ0KBKOF4EiolTYsqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqh5dTyF5Y9BDoCoFMPLfai8SJqkLs+k04K7Zo67q1kMyn1k4wbIBPzv/RH+ai4kudK
nNzpN9EOJaXo0KOc/9XEb09AHUqNPiKMXd6TmqYHnDE8EyhID5H/ht56af8vWeqFV3zAdArhq6j64Dh3Zh3Yk+tlQPW22L5SUWjdlWUY6VmR30qFNgPP8I7PTJJujGE7
2IxgPx4X0/eBdEw8eySRiJ5DxCzEkASNymFUZ4DxMUbNcm0jZkJUJy8xdjkHuDFNU0lOZQCOdtJ614qa720i3K53KcPSh2oTViOuKcinso44zrFTMakno2BgjqCmE9/K
yogm0Sa9h4GMq195YwJtiKpdTQe1P54xVOX2gkGNl9cbGBQfnvcKrUdPxCRA6TXP9Q9tSwhcCQX8a+HKNwZOZdX/xBbsQD/jjPOZLi8VNQpos9gr+qosvhbE3JhD8efN
3gRHoQ0bubQUMPVuAEVMOitPQgGgvhnT6E6HCAMb+XjlS0c8sH2LEVwanw9Sju5NnSLuL+gbYbIoYYUf18QzFYOooWm88MvOI7u8sMApOk9K5GAQ9xk1ZRdGxNbFTdoZ
9eAhsbYpcvuVPp86ImPIquWD7tHa5dDCubxNXUrXUd5aSRcoboxHyN6S+jbnPIay69zNUiOvbUD7bx1cmh+c1uSwAajdzqkui8gGD5m9o2XKiCbRJr2HgYyrX3ljAm2I
9rswH5Rl3UkeJz+f63rT75T9a/9FiYPrOt8HUEV+R81LF4omHtpUmYp6ePFaiTste8aglDVaJR29WmNJv6ePi69nQr2dgZcxiOyrULEE4I3KiCbRJr2HgYyrX3ljAm2I
bhPCaJgHQmhd4PWX/OFIGaxV2M4tpWvfNyZayXaI1pPcO/+RfPAiqwdk1+4exHDGnzdEbyQ46SXpqxEBFK7IjGZPUIaY8nnHEEtsz52et5eDcRdOfnzDCIY08vsxLu17
pAng4AbUtLk06d97+a0QbIDfPUfwK0M+0HHPtNLEe+IHtP/eXeK+kt+9Guoeo4lMrcN6J9wArhUYVhb/YO2VisqIJtEmvYeBjKtfeWMCbYiJr1+Y0WAaMj/ktP30L3Ua
mNg4vmkAlceraJi0nFyt2TzlKrF8k5nnIyBEOMqyUQQucE8tsKM4t/lbjxbOt2VH7Rurs7eq5Ev3eDKid+730cqIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mF
MWSI9gIcTJzNUvHq34GhZtWJr1Op3jRJdcUt3oDWbuDTfs6uZlgq7tih3U/vDEYC3MH3yNHRPOMmuAV3JC21M3IHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+R
mRM12/edwCO3mTJp9pC7fUi1xO8DYDrGVjgqpqt8unoXTn6/67T6oR+XnIxyC6UhlmJwqSxzcxgAuF0utn7RHn1IKEo2SdJnyzr0362qFc6ltknvXRHg2VsAKljpVOuo
sGwH78Sg+9egWGRNjKrEWxz7ocyWY6xBBQ2jUWsKP7QhnIqBvIRYhIsfo5+F1YKpyogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh2/uqxxiO0/E0uqL9u69w/r
1qdfheNm0WWcsL94VZ8xi2dvmCj1GpDUGUdC9XfTZe2m7YS3tubtxBs0tGrRWXq70yGRnPZE1s62DA8g752IHLnP5Pjl4sHgFuRC5wOFZuAF7Ftxvpc6QVBbtiw8lOj1
srh1QWjW5V0j+Ti0f12k3vHV9eWjj7OL0w+wUQAsJ9a2F8JTI8fckIfUO9H6EUKU6cdV+3ONhDnp7Kb9AzvcQnE/iLc0kxkagFkcIIvqNZWyclL/rs+tsr2Vlo2+g0Qj
hc4jSwzDsq2W8fvr8FGgKkGC5vWNn5PRieS6fTOGhFnKiCbRJr2HgYyrX3ljAm2IFdJkT329i7COnhM1KYxKodvQGo1kLX9Bh3H8ng+N6XciapC7PpNOCu2aOu6tZDMp
tiCa5ktzHlZh1e4kn7dkMpzc6TfRDiWl6NCjnP/VxG9PQB1KjT4ijF3ek5qmB5wxPBMoSA+R/4beemn/L1nqhUG6sd5iULngdjzVlxJ4fIvrZUD1tti+UlFo3ZVlGOlZ
PG6hVttv4VvUoq6tVVEUt9iMYD8eF9P3gXRMPHskkYieQ8QsxJAEjcphVGeA8TFG6XtqMe7KabpW0SvgxDBkW1NJTmUAjnbSeteKmu9tItyudynD0odqE1YjrinIp7KO
gkAgvdE+qSUXDmH0ii/idcqIJtEmvYeBjKtfeWMCbYiqXU0HtT+eMVTl9oJBjZfXXgmSDF62ETpmfL06qF4gePUPbUsIXAkF/GvhyjcGTmUMRKPyZYKcdiCuQAYuU0tB
aLPYK/qqLL4WxNyYQ/Hnzd4ER6ENG7m0FDD1bgBFTDorT0IBoL4Z0+hOhwgDG/l4DmqiLkTLwENuHv1yVBcyep0i7i/oG2GyKGGFH9fEMxXBw6Q19/mhgz5aC4kDmMfj
SuRgEPcZNWUXRsTWxU3aGfXgIbG2KXL7lT6fOiJjyKrXdiJ9Ub/MlTGg8VfX4FUCWkkXKG6MR8jekvo25zyGsuvczVIjr21A+28dXJofnNaUZUrVcj7C3bZBlZ1g46NK
yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+8mmDjVbNS4nMjWVSZwNDWQSxeKJh7aVJmKenjxWok7LXvGoJQ1WiUdvVpjSb+nj4vDWbgAxivmb6m9ATOKEDTb
yogm0Sa9h4GMq195YwJtiG4TwmiYB0JoXeD1l/zhSBlwRPKW6o5uOBCTHiZ6H/Nq3Dv/kXzwIqsHZNfuHsRwxi00rOmNDqPKQKn0VvS6wHFmT1CGmPJ5xxBLbM+dnreX
g3EXTn58wwiGNPL7MS7texteXZecWpYyl4LD+dHYsO6A3z1H8CtDPtBxz7TSxHviB7T/3l3ivpLfvRrqHqOJTA9XT6v07UFvQXkM4HwOt6nKiCbRJr2HgYyrX3ljAm2I
ia9fmNFgGjI/5LT99C91Gt+3ZnjheUdiBh/EpdxM7zI85SqxfJOZ5yMgRDjKslEELnBPLbCjOLf5W48WzrdlR/jzQ8vb6Yo+FUSH3HYX8mDKiCbRJr2HgYyrX3ljAm2I
bcx9A3euJafUPZh7l1vZhfCtfEgW6obuCTUEcZZmoVTVia9Tqd40SXXFLd6A1m7gZRRgRAy5QhYGcSNgWOauqtzB98jR0TzjJrgFdyQttTNyBy6pfPxUoXEONUlR82N2
BgFkoZbbTLQ27IEut7gPkWFmepDBG8CGogdhEWx1kyRItcTvA2A6xlY4KqarfLp6EU6ASyb9R9qZDOvebCsF/5ZicKksc3MYALhdLrZ+0R59SChKNknSZ8s69N+tqhXO
J+YrLZ64vkqAQqw9zGQexbBsB+/EoPvXoFhkTYyqxFsc+6HMlmOsQQUNo1FrCj+0tcQsxEl98CVnGfWUuTpRXcqIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKod
+DICnsPw8o80NPtZZXF3F9anX4XjZtFlnLC/eFWfMYvrftRSIhf558ahOXA9SdjRpu2Et7bm7cQbNLRq0Vl6u9MhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbg
zruiM6tLpgB19kYcfv7DtLK4dUFo1uVdI/k4tH9dpN5ubASDJP6LmHRw5J9w4uPRthfCUyPH3JCH1DvR+hFClOnHVftzjYQ56eym/QM73EL0qGxkWmeBv7jyDG1Aa5OE
snJS/67PrbK9lZaNvoNEI4XOI0sMw7KtlvH76/BRoCrOddvad2EkOdY6NUJYcijFyogm0Sa9h4GMq195YwJtiBXSZE99vYuwjp4TNSmMSqG6VDlY0LD4LjySPdAETZdi
ImqQuz6TTgrtmjrurWQzKYpHBAQYgCkX76hva5bMW6ac3Ok30Q4lpejQo5z/1cRvT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oVk2V1ZIMo1zTRcT9AL25PU
62VA9bbYvlJRaN2VZRjpWZYJcnBVnfNaBn9Mr/+eIPXYjGA/HhfT94F0TDx7JJGInkPELMSQBI3KYVRngPExRrHwjS11jDMghjjlSjt1gDlTSU5lAI520nrXiprvbSLc
rncpw9KHahNWI64pyKeyjoJmuJ5/aqVM2FV3xvtdoTfKiCbRJr2HgYyrX3ljAm2Iql1NB7U/njFU5faCQY2X16MWChUHetXz6p98lb5cL3P1D21LCFwJBfxr4co3Bk5l
LT5rOHI7w9Cy3EmzAKUdw2iz2Cv6qiy+FsTcmEPx583eBEehDRu5tBQw9W4ARUw6K09CAaC+GdPoTocIAxv5eCTYpl1Xnm7LMzqUYL6dqfudIu4v6BthsihhhR/XxDMV
h+Zs8oXqVMVqk8QhkV24xkrkYBD3GTVlF0bE1sVN2hn14CGxtily+5U+nzoiY8iqo2HE86iMMeFk+Y9ntPi5dFpJFyhujEfI3pL6Nuc8hrLr3M1SI69tQPtvHVyaH5zW
qslZMdlMXGIjgiKO8fMrS8qIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPvvL+0gS1a5RZeeAnlInqAo0sXiiYe2lSZinp48VqJOy17xqCUNVolHb1aY0m/p4+L
yHshRPE1KSdlVn+s6HcqUMqIJtEmvYeBjKtfeWMCbYhuE8JomAdCaF3g9Zf84UgZX4B4xk7bmJ1OgtLsCn9Lmdw7/5F88CKrB2TX7h7EcMYWBrtB7/o4xXp7/sPJRd5R
Zk9QhpjyeccQS2zPnZ63l4NxF05+fMMIhjTy+zEu7XvTJxh6kHsGuS4XFczWrAtbgN89R/ArQz7Qcc+00sR74ge0/95d4r6S370a6h6jiUyDTOckG0+xdEIPVYN3U0sk
yogm0Sa9h4GMq195YwJtiImvX5jRYBoyP+S0/fQvdRpca2mM1mhVeffIxWdG6YB/POUqsXyTmecjIEQ4yrJRBC5wTy2wozi3+VuPFs63ZUcrb0IiiwwzkVbLt1LquLA7
yogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YUR8llQXWlkolfzWwcq1Vet1YmvU6neNEl1xS3egNZu4Lc+t0JkdEfFZxMfh8fRXpPcwffI0dE84ya4BXckLbUz
cgcuqXz8VKFxDjVJUfNjdgYBZKGW20y0NuyBLre4D5FbVNF2beIC3EUyJg9W4nBQSLXE7wNgOsZWOCqmq3y6eiCBZ+IzGOGpFu8goixXBn+WYnCpLHNzGAC4XS62ftEe
fUgoSjZJ0mfLOvTfraoVzpmcHYwjz50n0bVx01C+1wCwbAfvxKD716BYZE2MqsRbHPuhzJZjrEEFDaNRawo/tJVFXFjW583ZK/BGGWhXqq/KiCbRJr2HgYyrX3ljAm2I
VOnKOtP+caPjsSiR3xSqHUSU1zeYjGDiVknWacsjE23Wp1+F42bRZZywv3hVnzGLTrf4k5F7jqYCBszRt2eYBabthLe25u3EGzS0atFZervTIZGc9kTWzrYMDyDvnYgc
uc/k+OXiweAW5ELnA4Vm4LCfet7VSdjsPn3mOfNrpzyyuHVBaNblXSP5OLR/XaTes4SF5NeWnpCfuADZiR/PS1P+ZXqkqj2Rjq/8l3cPYXDpx1X7c42EOenspv0DO9xC
5c3KdNm6MzmMD/cdZu+/LPTZsS7scfKgwlFwzGCf0RGFziNLDMOyrZbx++vwUaAqI097mIlRUEyHZ/mvyKnj1cqIJtEmvYeBjKtfeWMCbYgV0mRPfb2LsI6eEzUpjEqh
xtt4To3MoGf7U8iDidYymf8Sbv+7rF9B6egasVWcHjKwWip7t7P29mkuSC7gxY8kgN89R/ArQz7Qcc+00sR74k9AHUqNPiKMXd6TmqYHnDE8EyhID5H/ht56af8vWeqF
PFyM4vHgSMlxtYd9HE3q7utlQPW22L5SUWjdlWUY6VkGRCR5N6FYsB8kXEn4kRtEMuHGaFiqC0Va40HOdhiyS55DxCzEkASNymFUZ4DxMUbfvaLl77tyIMiSBZsHoIDF
KaJiHMDiUQaJQgKTBOvJka53KcPSh2oTViOuKcinso5ImKDGG/kbJktIviA+APuQyogm0Sa9h4GMq195YwJtiKpdTQe1P54xVOX2gkGNl9dB4QQ55NtACftF7YRf7P4U
+NYqKtNoL85OpJq2IDvczYuqgnz25efROE/VNMqcOxs2yKUInRm17Sfwi4NZWWjn3gRHoQ0bubQUMPVuAEVMOitPQgGgvhnT6E6HCAMb+Xh8oe4e/q3EksL+E/MWhIEa
nSLuL+gbYbIoYYUf18QzFRpS8/AVmEO6UYn6GMm6F0CnHqOgU55uXDWCN1Ydicbs9eAhsbYpcvuVPp86ImPIqtgKMk/KjmCNu7q8ZjaalnTOlJaKtLIITbM8GeKhPYmR
69zNUiOvbUD7bx1cmh+c1rc6rq90RTRJriVT2tAxFNCBtdaRBqeOTD5UUzy+4K+A9rswH5Rl3UkeJz+f63rT72iHclqaz/JkM0P1lpl/OCwJ1iKiFNUEULvk/WWTQ4G+
e8aglDVaJR29WmNJv6ePiwJF1DBQCnyLi4TGZEjUnqTKiCbRJr2HgYyrX3ljAm2IbhPCaJgHQmhd4PWX/OFIGfFHlZcjwt44k7g9ZseeLBncO/+RfPAiqwdk1+4exHDG
gF6y6gR2QR8DRhimIFlgDEd+8/x0979mmloRl34z6cCDcRdOfnzDCIY08vsxLu17CpheDRSbxitgDKeEi4csCITlfjm0JtbBwkeOXLm68fUHtP/eXeK+kt+9Guoeo4lM
I/TyMrQAY851TIuwbRqCFMqIJtEmvYeBjKtfeWMCbYiJr1+Y0WAaMj/ktP30L3Ua/LGMY9ba1/oTdB8okvEfBmVsH+Mvi+e/9LtMEveU2XIucE8tsKM4t/lbjxbOt2VH
6OXh9Y7F6S/PuQqd8im67MqIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mF0sayeN3UmbzbaiiYVp3Z9NWJr1Op3jRJdcUt3oDWbuCvnXZbsO/WQ5erieUffUTe
U0lOZQCOdtJ614qa720i3HIHLql8/FShcQ41SVHzY3YGAWShlttMtDbsgS63uA+RHv9xU6L83bM4iOiBJUoRGki1xO8DYDrGVjgqpqt8unrBxzedK8bhy1I6JIgq5ykt
vdDEE33/Y/o79/QXczL/aX1IKEo2SdJnyzr0362qFc5mrA0fzxv4XgytkpX89h0sk1FCxEbCHP5ya8GlIRi0/hz7ocyWY6xBBQ2jUWsKP7RyRXj0hXJTfnL9gkhiJQhl
bj3Ko4+CjH8yg9uuGxmZnVTpyjrT/nGj47Eokd8Uqh0r1CbVoEKw3CzlpbQS1hsKPUpsODFIrdbp1fwdkKAAvCsftTTX6n1dRRMNVJe0A+VaSRcoboxHyN6S+jbnPIay
0yGRnPZE1s62DA8g752IHLnP5Pjl4sHgFuRC5wOFZuBy7uB50uWrIKsliCCUjksesrh1QWjW5V0j+Ti0f12k3n0U3ppvrzO49isVRXPEHp9T/mV6pKo9kY6v/Jd3D2Fw
6cdV+3ONhDnp7Kb9AzvcQqXXZSm60XrfcB1KrebnegP02bEu7HHyoMJRcMxgn9ERhc4jSwzDsq2W8fvr8FGgKj1Kyb1wx4aySe88w34b1l3KiCbRJr2HgYyrX3ljAm2I
FdJkT329i7COnhM1KYxKoWRJmvG8T+dML3jWL7ytdlX/Em7/u6xfQenoGrFVnB4yO+0Mdd1lk+Gv/L0x7DB4GIDfPUfwK0M+0HHPtNLEe+JPQB1KjT4ijF3ek5qmB5wx
PBMoSA+R/4beemn/L1nqhf333RM5kUh7fML29tO+fojrZUD1tti+UlFo3ZVlGOlZgVfiraoxQFQL1TVl81jfRTLhxmhYqgtFWuNBznYYskueQ8QsxJAEjcphVGeA8TFG
xLbINJTlKrJh1Sshi7sitCmiYhzA4lEGiUICkwTryZGudynD0odqE1YjrinIp7KOegdn8uy/FnzDg16dIhZRMMqIJtEmvYeBjKtfeWMCbYiqXU0HtT+eMVTl9oJBjZfX
fe750UKuKU0KRfOTaBYM/fjWKirTaC/OTqSatiA73M2LqoJ89uXn0ThP1TTKnDsbySw2vN4tiU9b9W9uYbVdqt4ER6ENG7m0FDD1bgBFTDorT0IBoL4Z0+hOhwgDG/l4
1soQByiVJocjvuj4lNaug50i7i/oG2GyKGGFH9fEMxUxpwM0sDMhIuEXtLXHADjIpx6joFOeblw1gjdWHYnG7PXgIbG2KXL7lT6fOiJjyKq4bxDNeTwVcA/uWpQI0etR
zpSWirSyCE2zPBnioT2JkevczVIjr21A+28dXJofnNZIvVkwxVV2rmTpLKElcodzgbXWkQanjkw+VFM8vuCvgPa7MB+UZd1JHic/n+t60+/Qz2PNQDmZ72XELSw9VA8x
ayn5XBJoVZRbANEMi+NKfJnlbEAOZQIDJXV2A/etOu7KiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiKoGj5MN2FrbDQGGH6xddEs3c5wuSWL0U3fW+ed3JyVW
g7/lw4e3tjxkHreCiucDFgP81xEf/yCOtXCmcu1t9K7KiCbRJr2HgYyrX3ljAm2Ifshma5gZ3m5WUZsPRTH015MEygrQ9+FtWyjlwNGLxA+vV2yXOtafyQM1aErUfdNv
5mC6Z3xj/Cp09clXOt/rzPdzNf6fpzF8d3g+zBkXxjjKiCbRJr2HgYyrX3ljAm2IxARU36a2APFypw3tFicy+85ZQBPss/TvsyZ9tRUY6mWLYGtvY/Vs1h2pytLRB97E
gRrInBgZD19HN9j5BZzno7irG3IRRCRrU8dALofRyyjYjGA/HhfT94F0TDx7JJGIuoiCPzzT5h7g3UlNEM4jRLa5PSTWwNdSYmQla1BUWQ7KiCbRJr2HgYyrX3ljAm2I
NmWWg12F12lg4BpNV1U8x5XR6mMzBmkKbiuqARCX6+dBJmlIU7ajV4C6nYrYNjCXKMyNAvbEdOTszf2KQxnqJcHO3OxcfH/rOWex2vgsLmckF9dvoI2mAgTUeUHLCVdI
0yGRnPZE1s62DA8g752IHPj97RxDFrjr4QcDBRgAwW3JkTx38zJquLieRZiUlINhJnZr5EurXoMNQst3AxzL3tE/XLE7d/FK6qJ1ErpwIEdIHqOfEHsLTpHSbi5HZyKy
cmNCpBnjWbsQW9+auUYlAYzyRSy5917B74acfhXx+g1CDY6kpPPo85HB198p+T1VPWzu1WVz94cYTu3XYoQ+FYei8NYwyXkZeggI56UPn5MVdhHqbZnppnRnAP6kv77c
NJcVnl8nC2lJnazY7jtP2VBXDKzdsLlbUmJ6AgiVKLzROigIFlib0B49QuLx3JP070u6lR7N0aj5AzJlvr74/B6woIt5DBGqFg2eldIFnPByKYVyefT+bTR0DEfJNVrh
/1H7o56cXQFh8dCv4RWT3o71D8iCvw5rfsys96cMKvoTfCYuxJR8xqvwWlS/F3glW6Y+x6+dz/xqtGqKzGakffaHQKAYawCYqvWBU9D32n5UJ85ITb6XO/AvolOAW1aY
KnIMB9KcfZHV+WmAiMOGQUd0IwgHnfu8CDR2pJUv47qYk88PUh9xEvGxqQDYhF01aYTXYsfI0OkB7OPO+5ZOyD4gfLIz5h0+K0oXuKhg9TTuRoz1bKvhMx02vJAveNPw
I6MZOJ+JU7iLo+xdUSBlEogkScrPGn2suDPtYWT77jodtuf3RZZL9mfcmDDMlUTnsECBbdgdd4Jyfk9VZ2LW+JL2n9mrqUsRfDW1LbmctW2NPhyyZTl3krzf8rJ2bF/P
7xNsfSnawPp0418jdqIPWHzjPVpKFYWvK0ep2ykku4CdXnUNvkNIyZpSu+LHQf6xoG+TQl9IdvyJhuLcwZZtgOXN2D8F0byLJ4Akjo1vFWOmmx5t+tfsJkmoTIPWyOrF
jEsF9BOsBJdta54FyZvg8GtZ5g5m7JuWVuKa0LNnibXlgAPpvBFpCOFgFuFFix42/fA7wzRFnddyYkIr5iMzicqIJtEmvYeBjKtfeWMCbYgupPBtmBhLIFiVKVFXC1bM
SJhpOFU3JEBDrxHqs9QEr8qIJtEmvYeBjKtfeWMCbYhAyaqwkAgzq4ApJkwTRqQMRG1bZxaWY7/B685bBDfEMMqIJtEmvYeBjKtfeWMCbYiOEeq51Jn2VxuzCmHvwpvo
pv16ffHTEUlC9z1UgLaKHHDvRSfVD0hRzob3Uax5dcCgU3uAd5P5mx4yFH6qOu0ikJyuNncdtmCmjwEFnh3GAy5ikYiNpSLu1/ezzjFq4+vU3MAjvbQ+ppjF4yhvqEIt
BbcYMLGxFf7jqt5GR2XSMsqIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17Y1Bt1tmsdKFYAiXn0R565zpvG7Rq1BIm++JChRdCpTNqomAJPclZBfWv/JSelZJ3
Xy1Y/SKucmbXSi6EF1hbYD1vJ5kUtYHPkyI525LqSgVPQB1KjT4ijF3ek5qmB5wxusOZ03wk+7zv6S9F4R/iDeSlV3P8KTsnpYOsGxat/XapBA58fpzmVa3b7qxbraMI
IcsIPWnSZnuVsm6Mtakl4HFTQ0gcvXqvk1d7T2wkurfKiCbRJr2HgYyrX3ljAm2IEx4urYUoEPuelpFBu9pbHpFVWpNmXmFe12IGwtYAfoCUVNyq2AQPD9kvJB4JjOsp
ziejpzfwHt54yBEEAOsU+8jmVqbhS9+ygCg4xSkZSJS90MQTff9j+jv39BdzMv9pql1NB7U/njFU5faCQY2X196nfnAN8ZIUagrOgjMzk9pWapOQ5OY7MWfmsHTheYcS
CwwAcvtg7iYlCwF42KyIGtZRfECrAsIHbKJE9kogjTAvXzKHvex7mvt+AdjW/17PfUgoSjZJ0mfLOvTfraoVzpadnmUUF9tCzXGoZ+EtNU/KiCbRJr2HgYyrX3ljAm2I
YNLYKxdBjjxtb6GvKOUTFIiTzaeBQzdz2bF8pd5cNDLKiCbRJr2HgYyrX3ljAm2I9eAhsbYpcvuVPp86ImPIqpNPkJ7gD/XGUjX5N6qz8Ve+Rgtf+aIwriJGmjgpJ6RX
rsiVPgYhD1stOQGflq+3eDdznC5JYvRTd9b553cnJVbKiCbRJr2HgYyrX3ljAm2INFiVMTvyeS7+I3Z0qRQ0X3igFh0Ld6lpUrixOWI1RGvOu8Yukwrzv9xXwxo54ngL
cJzhsIlxNnjOPUoTg6WZxKxhqrW/8yzz07lMxb57St08rQ/H+Chw6MmitXJ91FsC7P7kec8cXWBcdxverVThJkmV3UcDeLGhA/7PNcP63UwvvmNDby730bqDNdanrDVn
hdGjW52EIvIfw2vdC99BIMqIJtEmvYeBjKtfeWMCbYhU6co60/5xo+OxKJHfFKodqQNZ1U/+TLtpQRQHXuDh68qIJtEmvYeBjKtfeWMCbYidohm+coC6C/i9PN9CtkEn
L3GqXvCz7yJicpPflpna0DLhxmhYqgtFWuNBznYYskuJr1+Y0WAaMj/ktP30L3UaounTuyZsuHX0waCszGX6vkCN/ND3XZvaB8pjXVLWrgP2h0CgGGsAmKr1gVPQ99p+
STjFH+mb/MbkfV5ZW3hf20EmaUhTtqNXgLqditg2MJf14CGxtily+5U+nzoiY8iqq4l8Nfy0dN2OU3UzdeFDIcmRPHfzMmq4uJ5FmJSUg2E9DaBNeTZ/4lDYiGiRR45S
2UJXRRp9SFHMzhyE40MUMJcBk8UmWwf7r4JmpLeJJ9H0RERiZUup8QKDSg8ekRnZeZeLRwEE3MinVTuLvmGoII+eCHvSOgNhLtY5UadribDY1icoU1jnFOVf6U+RDgl9
L75jQ28u99G6gzXWp6w1Z+8TbH0p2sD6dONfI3aiD1hffjDKjWFZ2z1UMFrVfr4KVOnKOtP+caPjsSiR3xSqHQxho2El/5iYVGXTBT8GY9bLxKHBtsvT1ljtQATxvRZK
YrVu/YCaUWSjIu+r1S9bcxV2EeptmemmdGcA/qS/vtxbFKQbHLttSxZStTV9w5liAFBbDviLnpbjJVFgIhg7z7GrRPOxL1ZZhnKhdbvXb4brW++djTHn//7SO2s2Y9Ye
9odAoBhrAJiq9YFT0Pfafs75ZK4RrN0XbAjOBuhrJRSjXf5M6pxUJaD6whEODKMCRP5WgZpjjT10r/GxJyAbAauJfDX8tHTdjlN1M3XhQyHhsgeBRaLW5blz0nv6+dao
KMyNAvbEdOTszf2KQxnqJdlCV0UafUhRzM4chONDFDCXGEFER09NLos2DtV4QrWkgp5po1mxHS1QsNMZxrFTQ3mXi0cBBNzIp1U7i75hqCBz1Q8E11WdlsXwE+UXlyhU
0nsdEcKwtwiQqWAQlwCO2y++Y0NvLvfRuoM11qesNWfvE2x9KdrA+nTjXyN2og9YCGvHj4Wd3pJCyiFvJp8141TpyjrT/nGj47Eokd8Uqh0MYaNhJf+YmFRl0wU/BmPW
2bPoOpfcTwbFb0FbraCaimK1bv2AmlFkoyLvq9UvW3MVdhHqbZnppnRnAP6kv77c071Ryi+qiA0Hhdug1eNnNimwFpr7r3fIpVdYnA1fXcuKyKR3wFwIHeHPCGzekGAL
UxoQeWydCxDIplUUgtQSr/aHQKAYawCYqvWBU9D32n46ZVAyd2auanP3mbakox0S2nwprEjEJ/BEkk9longSKTZlloNdhddpYOAaTVdVPMeWsb+5A6B/yQCHmCiI0hqg
AnmZQIT1L+hYD9RcIrxTlyjMjQL2xHTk7M39ikMZ6iVwgRPDf/0MIt4IukV59bRU1A6Y4zXqsfGOQk9PLoLFvU9AHUqNPiKMXd6TmqYHnDF5l4tHAQTcyKdVO4u+Yagg
+NYPBzWB0/peGzXXO0GwIUmV3UcDeLGhA/7PNcP63UxU7uqJ67LifigoZFSOHHoezFzDhyoiuQCyF3vnaXB92cqIJtEmvYeBjKtfeWMCbYgefHETnzHurOyvbf954PnK
N6508f2x6uWGDBzyv5mPO5d+4MgSYTCU5FJ+KYWwOd+dohm+coC6C/i9PN9CtkEnmLOfZnkO+S/ykdbs1PN4lT1vJ5kUtYHPkyI525LqSgWJr1+Y0WAaMj/ktP30L3Ua
AlXD5PZIK6ZGaYnecb65smAMhM7uGrm8FzWxlTypAgz2h0CgGGsAmKr1gVPQ99p+OmVQMndmrmpz95m2pKMdEoCmNxzirTYd7fXcs4sXVIQ2ZZaDXYXXaWDgGk1XVTzH
lrG/uQOgf8kAh5goiNIaoHztZ8/w1UxPq3rwUrUlxDsozI0C9sR05OzN/YpDGeol9MEKdMY7SA4RaXT5dX+JqddPiiF7BWEzhum9Grrdmrcp4OTXOviXMTHM29B1LqGF
PBMoSA+R/4beemn/L1nqhfwGOhJxbGluJB/ixWNM/4ujJ2f/BWdlPrqav0zEHAWSVO7qieuy4n4oKGRUjhx6HtxNVTyrJcJJNJwB/K0ICjVWapOQ5OY7MWfmsHTheYcS
HnxxE58x7qzsr23/eeD5yl5/vxI/XqEmevWJotB2YdfKiCbRJr2HgYyrX3ljAm2InaIZvnKAugv4vTzfQrZBJ40/HQ7wkqQfC7ylxxFTbRn7rICpy6vrQuFpgCGDT3b1
ia9fmNFgGjI/5LT99C91Grr3RGfH5m6DjGDLnXSMUDqxUpBEHIYNAgisGtBZb5zqFKAcqMzyyv4GnLnBTjZMqZcF8kgtrSst9snoJVzHFj/KiCbRJr2HgYyrX3ljAm2I
9eAhsbYpcvuVPp86ImPIqiv7Z5piUGdNYHFs6eY1Y70hvBPv4szoA2bQnE+kmNvEKMyNAvbEdOTszf2KQxnqJcHO3OxcfH/rOWex2vgsLmckF9dvoI2mAgTUeUHLCVdI
T0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oU2uc5g2Oe1H/56WEnpENnZjlk1bDAmGXGBgFyCOlZONVTu6onrsuJ+KChkVI4ceh7T/QlWbTbsaIHkcd/f7edx
M+rZT0ajHz7sixcQqGUHAx58cROfMe6s7K9t/3ng+cqY0NLYrjQKfbM6fXVP5fElN6XC52fW5cz7b62pCMp2A52iGb5ygLoL+L0830K2QSf2/1P6K3V8Vev77Crkg5vj
p96W3VtnIC3fvWoipO87QomvX5jRYBoyP+S0/fQvdRqpI19qwryT2npYg2oNkgZFbDDESQ65KZV9eEzUwDjSi/aHQKAYawCYqvWBU9D32n5UJ85ITb6XO/AvolOAW1aY
rhZWkKIENaTfNEejVTmrpkQqK7WYKpM5gdYPN+TU+Mcr+2eaYlBnTWBxbOnmNWO94oya9w9tWvW4KHP8ZKPv8k6nVIGjeVcKFzZ5nxOWub7BztzsXHx/6zlnsdr4LC5n
7RJb/9kOnvUS7RTAWpVh1Cp6EhbEeGiej4l4/uPrgfA8EyhID5H/ht56af8vWeqFOTl5MsSDYY2mE1Qj6KVvb/Kn/adPWLa9Q7nimM2wms5U7uqJ67LifigoZFSOHHoe
0/0JVm027GiB5HHf3+3ncQE6Uxivj/kNWWHWaRIwaJsefHETnzHurOyvbf954PnKmNDS2K40Cn2zOn11T+XxJab4/aEWeU195TUVMHbq8ACdohm+coC6C/i9PN9CtkEn
9v9T+it1fFXr++wq5IOb4zQvUjofpDUJgi/8EpXEmSKJr1+Y0WAaMj/ktP30L3UaqSNfasK8k9p6WINqDZIGRcZYsRGgBt5FiwE6FcJmjRv2h0CgGGsAmKr1gVPQ99p+
VCfOSE2+lzvwL6JTgFtWmA7f6diZ6LcPrbzrI1dj4T08pxx28HdEtnWGBBNlsv5wgB9qsfweS9slr1Le8fyWWtFYpKpzkRf6HRt3vA2syGcozI0C9sR05OzN/YpDGeol
KJJn56XQC6v8BkzbXdxv8k1/dFQI+bNoTdA3CtXKYvRPQB1KjT4ijF3ek5qmB5wxeZeLRwEE3MinVTuLvmGoIHS9GEclc0w38oV9nQyi2dNJld1HA3ixoQP+zzXD+t1M
VO7qieuy4n4oKGRUjhx6Hh0QS1w27BxVTyOEBXPW+DDKiCbRJr2HgYyrX3ljAm2IHnxxE58x7qzsr23/eeD5ykBxz2q0IpuGpDrAlwne1iPKiCbRJr2HgYyrX3ljAm2I
LqTwbZgYSyBYlSlRVwtWzDCPESMbaD+NVaJYQWhGtCTKiCbRJr2HgYyrX3ljAm2IKbAWmvuvd8ilV1icDV9dy9pBRWzWa4tXEhuAFOTUEI6XsKCD56b+d8pLuPYEFPcW
FKAcqMzyyv4GnLnBTjZMqcxQxUmeV29HP1gqX4rRAvtyY0KkGeNZuxBb35q5RiUB9eAhsbYpcvuVPp86ImPIqoAfarH8HkvbJa9S3vH8llpqBR17tWQpht24Vd8GxHAh
PQ2gTXk2f+JQ2IhokUeOUrRdI47NwujMT+Ti30OJEglUTxQ2Dc2SQezl5vSWbXP2T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCAgdAy8kJ8fiE1xMrYpTQkO
8qf9p09Ytr1DueKYzbCaziHLCD1p0mZ7lbJujLWpJeCoO47DyXYZ/rK/4lGYa3iGMs6Yp83sbEijSPVFltsRMFTpyjrT/nGj47Eokd8Uqh256UAhN3bv55NfzSmuKp4a
2bPoOpfcTwbFb0FbraCaii6k8G2YGEsgWJUpUVcLVsyqmapYp0n3Eoifipi6/AlsFT+c9sG3BSRt7uxphnHYzCmwFpr7r3fIpVdYnA1fXcuykd3BWaN5sul/4djlzOLj
yogm0Sa9h4GMq195YwJtiOsuWmbEdf58c7NWvSnS7BfKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKqTT5Ce4A/1xlI1+Teqs/FX
vkYLX/miMK4iRpo4KSekV67IlT4GIQ9bLTkBn5avt3g3c5wuSWL0U3fW+ed3JyVWyogm0Sa9h4GMq195YwJtiNG7N7soTyV31eElYIiZuMiRD8PBjEBPPcILu+2mTiuJ
XsMo/Wrb1ululL73jDmbzhZ8YboDvNJhIJyuVJ7OG5LKC07R151eAfqW9XTIMT9RoGqbrHTFDMVdbHO2n1tV8cqIJtEmvYeBjKtfeWMCbYidwFtoK9RltnRHcF4zvllK
9QG9FuxxgYlNMGmWzzyRfciGEPvq+Z03vanUQJWE3b3TIZGc9kTWzrYMDyDvnYgc80s1u2OqHYTm0Fd/2Mp/6KWRnKhK+FRF8UcAIoQlSvDKiCbRJr2HgYyrX3ljAm2I
i6R+zFDVDArB+R50NlHD2X2aOHn+u9yUV8hBGw/VZmoy4cZoWKoLRVrjQc52GLJLNmWWg12F12lg4BpNV1U8x6uJfDX8tHTdjlN1M3XhQyEhvBPv4szoA2bQnE+kmNvE
wdqysPuD8M36TcA/bSQFwYYYVXZDH0M1DIKKRVIx/EqwhlnUgcagkchph+haSJPmQSZpSFO2o1eAup2K2DYwl4EayJwYGQ9fRzfY+QWc56OjaqOmB8Gbu+bzvDlR+Fdz
yhv2DAx6htG2rwiEmWl+ZRSNyUk5VeZ7+SqbWWfc3KKAXbtaWIS3elSY6NpdD7PbW4t+El3yqAzVo6Ueev9Q7lw1M60Jz4ZwSjJZd3axuO7S9n8LkPi7FXyEZHTrIDFz
SgEQuSBNhFMpCWNGJR8ChVRPFDYNzZJB7OXm9JZtc/Yq8Cd9J+SlOu+xBuUPyZ3cwca5JFkF5DVCXFh2+PcTmNP9CVZtNuxogeRx39/t53HC8k90SngXIPuXw2mGsBfE
bcx9A3euJafUPZh7l1vZhcu6bpf0koypEhaaTKQKyZx0qZQRJ8MER6fNGs33p4qT36XbMRKQePRpdT6uwSSooRT5woCDkTCoNf17S+G9NfHIUp4yrsrkjJK4f9NGSXWb
h6MIrFFNlIyHnfqIq6FaTHmXi0cBBNzIp1U7i75hqCC2DM8PyXpUDsCmHtD3SKfj6rSQdmbmu3bjd8udEHqQslDHbpfe1euVF6ljsJs4EeIMV7GKYfAi6dtC+Zgv/uO4
n/klliVLMhZ5RiAytKoqtCfsjfqSE7BuOQ8I1493hLJUguCL2m2vpjJ2bKzelzzAlxhBREdPTS6LNg7VeEK1pJERLsC1IlWRGd1c2zLeDPbbskS6rZvAxa5+jrBBT3uc
60yrTofVOMuG3l7phW6jb6g7jsPJdhn+sr/iUZhreIZmgmpNWLWJVEUhiZ2nvig0esvYt9Cvezix4fT99y7vJWVQ+qZyzRo1bKnidehPSnWSyv7mlCuiNFcSWG5SSuJg
VovpwjX66oeTMs7V+XIbqPb/U/ordXxV6/vsKuSDm+M0L1I6H6Q1CYIv/BKVxJki9rswH5Rl3UkeJz+f63rT77111QhUeY0Vt/OTOatyTvPSQ43EBgKroxSYDs3ORJtM
2/ZlQsl+mDj7nALuZBsrJyzF9A/TKeFm9mRiN8kYid6MSwX0E6wEl21rngXJm+Dwa1nmDmbsm5ZW4prQs2eJtVTpyjrT/nGj47Eokd8Uqh3NLVrjjTimRkzz3aUR8npK
yogm0Sa9h4GMq195YwJtiKwP4yzBr5hlTX1UqpExRu/qvxYGoHGCuAX02EgKolLI0VikqnORF/odG3e8DazIZ94ER6ENG7m0FDD1bgBFTDorT0IBoL4Z0+hOhwgDG/l4
i5Wv1fNdOT8nROu0jTK4xsqIJtEmvYeBjKtfeWMCbYh2N3LuDhJ2CYsCxCyFfBcOnbwEU8aQLSrK1q2/DdHA69N4D+wHk19YOJEoBAac+tVyBy6pfPxUoXEONUlR82N2
RPSVlqBUKpiz/b3JoD4gIDCPESMbaD+NVaJYQWhGtCRJld1HA3ixoQP+zzXD+t1M5aNrQml3xR4iCFSUilJcEUqw1tfc/JnebmGSw6rUkdTKiCbRJr2HgYyrX3ljAm2I
oY4ZFtMWUeI69RCmMkyCzduiCEtzO7rbXQFoyKp7YuVkSSWOK5OyJ0f3cKOFeykQQsdjCaTmfg/wrR+cdLwJGa1VmbHBSA/7PYqURZ0Xpy7cTVU8qyXCSTScAfytCAo1
M+rZT0ajHz7sixcQqGUHA4mvX5jRYBoyP+S0/fQvdRoCVcPk9kgrpkZpid5xvrmyYAyEzu4aubwXNbGVPKkCDN3YIZnCtcfZgKOTAI+c6sy0KLnfOySySJ+1yrX5vGKc
tz0+H6Kata5ZKVpZsETs8AQkgHhgJpwSdmaWWp3h244V0mRPfb2LsI6eEzUpjEqh2Z4h3MDRCDEjtBXMW2w3cIOP3CrxBZ0DXWDdD8DV+je9XyBoyERARDr84jKP6d5S
cgH2jt6MUonEdizqHQ7KNMjmVqbhS9+ygCg4xSkZSJS90MQTff9j+jv39BdzMv9pbhPCaJgHQmhd4PWX/OFIGb8XtI+WPTRB8Qb2/KT+nT4CD+Ub2TcuiMyZVl6wfe9+
ncBbaCvUZbZ0R3BeM75ZSiDGL5Q71auz8mEhd97buIndnFF/pAXdg6FdAIyt1HS9l2WpShs+i72ymkJnoXpJqpI3DT1waeDxQLTO5qtyfNVDdEBUH1fBr0YhhKlapneS
yogm0Sa9h4GMq195YwJtiIukfsxQ1QwKwfkedDZRw9lQgMzrB1mOhS75DpAbMvYDRdy5PvRglrwdSL+aTHC2TTZlloNdhddpYOAaTVdVPMf1t4TqmF+DK87kmRSb1Cnq
R37z/HT3v2aaWhGXfjPpwMHasrD7g/DN+k3AP20kBcFDLf1xBEmw2fsUr3K5S/91sGk+m0gqMN5GZlv3RTDGQMqIJtEmvYeBjKtfeWMCbYh9SChKNknSZ8s69N+tqhXO
AQYEynmDGqiWzOhuYMT7ZKVjCWUq1lGm2UiZV2CVqsUUjclJOVXme/kqm1ln3NyiV3PFNLVwGqZHwu1C64l0QmSn9dj8yXDYuRCxZEqyw6nKiCbRJr2HgYyrX3ljAm2I
ql1NB7U/njFU5faCQY2X12+ZjXM8depxJx5+z7c40DrKiCbRJr2HgYyrX3ljAm2IVAQrHhRdPhBfekpiq7q3cm0RGbwsqUcnRm0WTJz/+0HKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YVaOAkKg8t6xNKZo2Hm+9WLyogm0Sa9h4GMq195YwJtiN+l2zESkHj0aXU+rsEkqKFZvA0dgM4HZ6bYEdFYpjle
dG8cFsWcVMfy3KpdNwWSCE9AHUqNPiKMXd6TmqYHnDE8EyhID5H/ht56af8vWeqFkFPKzbyzKeOzRUhANUHQVMqIJtEmvYeBjKtfeWMCbYhQx26X3tXrlRepY7CbOBHi
FbwZ8b487l+04dnCuDJqor3QxBN9/2P6O/f0F3My/2mDcRdOfnzDCIY08vsxLu17tpOsZz8YKYkExTeR391K8M58t7JkjdkM7RVfTU/w39qeLF+C2KCgIOFSqtYkwROa
uwOPQ25eSAg3nYe6T2QWQX5hg0AT71nXvZyEBSVZkZfKiCbRJr2HgYyrX3ljAm2IoFN7gHeT+ZseMhR+qjrtIhg6yJBvXwNcMct88BdG7UWy+U7twSdIO7DGbdUaIUjX
9Q9tSwhcCQX8a+HKNwZOZYdYtHmlcEiCTQbMMWSDf7NZn4UANi/OXjUMqi2Igy8dyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+/Qz2PNQDmZ72XELSw9VA8x
yogm0Sa9h4GMq195YwJtiGDS2CsXQY48bW+hryjlExSIk82ngUM3c9mxfKXeXDQyyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhZKODriqAGJStbrevKmGRQ
ho4Bk3CGftO55JtjjGCmgMqIJtEmvYeBjKtfeWMCbYjERtfOPf03lhTZXmjLajDFvkYLX/miMK4iRpo4KSekV8qIJtEmvYeBjKtfeWMCbYjeBEehDRu5tBQw9W4ARUw6
DfnOIPsucGXhpFwNkbNeg5ChsDW+564t8Pfdsn8uBQN+djVNu6+r+RCAMbghsxOlzxC21xL8hfi5fFELwA9qPqF1w1GnpogKGlcsiPyuVnLIhhD76vmdN72p1ECVhN29
yogm0Sa9h4GMq195YwJtiM/pZPEZhq3IXCT/N8ri7nNLYOI+uNojXevQ9oT40D3n3fdyYNKT1Io2V6H63wgKoU9AHUqNPiKMXd6TmqYHnDF5l4tHAQTcyKdVO4u+Yagg
cSgMgEYwnThNilSoK9BexcqIJtEmvYeBjKtfeWMCbYhQx26X3tXrlRepY7CbOBHiit4rokOpaizL2A0yyKuQQ31mwD3CEYtXA4GZ7WwI/NDeBEehDRu5tBQw9W4ARUw6
K09CAaC+GdPoTocIAxv5eNf7febNJq867oHjb4s7nxnKiCbRJr2HgYyrX3ljAm2Idjdy7g4SdgmLAsQshXwXDqLP9PpOTtbjM66jfhhF94ohvBPv4szoA2bQnE+kmNvE
yogm0Sa9h4GMq195YwJtiEVO3OPgHLKAqfJChKsasjL31lT0h3gqRiP6OdFLVZypcmNCpBnjWbsQW9+auUYlAZ3AW2gr1GW2dEdwXjO+WUppWkNIkR52+B1lg04MPUyh
lwGTxSZbB/uvgmakt4kn0Uy/4VG4PBZLfml+3MRz7RptzH0Dd64lp9Q9mHuXW9mFy7pul/SSjKkSFppMpArJnMLyT3RKeBcg+5fDaYawF8TfpdsxEpB49Gl1Pq7BJKih
cicZweWlvEswe9VnG4WWa3wBsaKbAXC+3OGiD5pfLhpMGCTfHWX/c70MsyNHTs8nVOnKOtP+caPjsSiR3xSqHQxho2El/5iYVGXTBT8GY9bLxKHBtsvT1ljtQATxvRZK
rA/jLMGvmGVNfVSqkTFG73f0RJdOcYZLMskPYm+HrsVLbYTiCDt8iUfqA2gWgnQyJ9nKa7jaGYmf2oQ3GbMFvHRDKVZNP4lSwf13PICjvgMzlCveq0vMQePGY8kWctn/
W6Y+x6+dz/xqtGqKzGakfb1fIGjIREBEOvziMo/p3lK1Y53WfeyvQIvtQZD83MrozGZZcwqk2Oss/hzzCBUyKCtygoBgT92SUC0K1xHsm9rS9n8LkPi7FXyEZHTrIDFz
SgEQuSBNhFMpCWNGJR8ChXlKRnv87KxhwcJZmKMxBt4q8Cd9J+SlOu+xBuUPyZ3cBHQeEgmFpU2V2oZrW8ortO8TbH0p2sD6dONfI3aiD1jfhUTn14E4eQKv0bVgGJYm
9rswH5Rl3UkeJz+f63rT77111QhUeY0Vt/OTOatyTvM0c2Oy0SK3yVyui5fTmWe72/ZlQsl+mDj7nALuZBsrJ/g9B4LRSs33D6Zx4I6x4TBIHqOfEHsLTpHSbi5HZyKy
dbPar8C6vviN/hvkd68BbimwFpr7r3fIpVdYnA1fXcuxq0TzsS9WWYZyoXW712+GxlixEaAG3kWLAToVwmaNG93YIZnCtcfZgKOTAI+c6syCArVGlwEyH9dSs2GwGuOd
0/0JVm027GiB5HHf3+3ncVZqk5Dk5jsxZ+awdOF5hxKBGsicGBkPX0c32PkFnOej0XXXLgbpccufiV0/Efn0uotga29j9WzWHanK0tEH3sQUjclJOVXme/kqm1ln3Nyi
gF27WliEt3pUmOjaXQ+z21G3ry3KrXHlQGCTBRJ+qs1Nf3RUCPmzaE3QNwrVymL06cdV+3ONhDnp7Kb9AzvcQjv2I/ihpPDXreHM7jq5yxtw70Un1Q9IUc6G91GseXXA
ksr+5pQrojRXElhuUkriYHn2nMmMJoOkHYsMsd9Tsfl3plvj0+DwgM+qrgBr9My3yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUbboghLczu6210BaMiqe2Ll
1yeKbPAQ7QYSbInpH7pkkkLHYwmk5n4P8K0fnHS8CRnhB4i7RFNp7oT7X0hIxZQLaxP3IZci3k0TRBAAwx3vUkCN/ND3XZvaB8pjXVLWrgM2ZZaDXYXXaWDgGk1XVTzH
lrG/uQOgf8kAh5goiNIaoAbZhRxQk/b115uvDVp8fYu9JUi1COi/uBgiJFQM5xWDhhhVdkMfQzUMgopFUjH8Sgdx+yzjydMPbtzud3JeWvnKG/YMDHqG0bavCISZaX5l
g3EXTn58wwiGNPL7MS7te3wuCEegFy4Sxost61XiCXTkpVdz/Ck7J6WDrBsWrf12I59VM4+Y2FuID/yHDipKEduyRLqtm8DFrn6OsEFPe5z17ET+DYV03lMnauL4fHAO
cVNDSBy9eq+TV3tPbCS6t3IHLql8/FShcQ41SVHzY3ahjbooTTPfJWrbBnqAdmZMA/1sSabum0a5+IQ7CMWTSqjyXz+U8VmzgJ9hwCIq/GgfgOjlds/lBEgdFn/gEv45
OmVQMndmrmpz95m2pKMdErYd7fKrWDa70kDmD7Hkv7LoYZX65StPHIV97J2Z3qTb/Q3CNWg9Cly6qTkokiDXWGEW8yNkAhhGNQ/qptpaKglQSxrg7f6n4Jn75yG8WZrQ
z+lk8RmGrchcJP83yuLuc5K6nMR4mHSYUGkTpQpzg0qpke42a8avDa8r8kKYOYu9rvuz8E8rXcqHJVE8bbEOFzwTKEgPkf+G3npp/y9Z6oVHwzRbPv3tGRCq5ap36hE1
yogm0Sa9h4GMq195YwJtiFDHbpfe1euVF6ljsJs4EeIMV7GKYfAi6dtC+Zgv/uO41wfFMPJFsyStJ9zq/W/Qxd4ER6ENG7m0FDD1bgBFTDorT0IBoL4Z0+hOhwgDG/l4
cw2+qOIWbvji8bh1lQa4BsqIJtEmvYeBjKtfeWMCbYh2N3LuDhJ2CYsCxCyFfBcORAY6+bKXhVHR8NxH6YHeiHI73gMzvv+1OfGMEuyVGhfKiCbRJr2HgYyrX3ljAm2I
RU7c4+AcsoCp8kKEqxqyMqcbox/OBuGs38fpiSJJYwTKiCbRJr2HgYyrX3ljAm2IncBbaCvUZbZ0R3BeM75ZSvUBvRbscYGJTTBpls88kX0kF9dvoI2mAgTUeUHLCVdI
yogm0Sa9h4GMq195YwJtiBJGqJWn1t/qGroimMFAGFbbmNjAg1IYfBpCGrbKiFQkM+rZT0ajHz7sixcQqGUHA9+l2zESkHj0aXU+rsEkqKEU+cKAg5EwqDX9e0vhvTXx
NrnOYNjntR/+elhJ6RDZ2UTogJKXOvj2i9jswBX8gR0efHETnzHurOyvbf954PnKmNDS2K40Cn2zOn11T+XxJTelwudn1uXM+2+tqQjKdgOsD+Mswa+YZU19VKqRMUbv
AkbjYk+qcfKO+1ehMddPWe8TbH0p2sD6dONfI3aiD1hffjDKjWFZ2z1UMFrVfr4KFdJkT329i7COnhM1KYxKoSEtpyJzxUvTubbO+dNMWvpEd1pM2JHvTr7hEV8ZJt9v
vV8gaMhEQEQ6/OIyj+neUh987aLTnUqU5WBDSxbwAsdIHqOfEHsLTpHSbi5HZyKyve0CGTjPekXxy3s/speLwqpdTQe1P54xVOX2gkGNl9cJjDpF6GKRKlYydR5vn+/g
lZI1zb/3WoHNywl6uq4IuCrwJ30n5KU677EG5Q/JndzBxrkkWQXkNUJcWHb49xOY0/0JVm027GiB5HHf3+3ncW3xa4I8yqsJjwjV2j9MZzhAyaqwkAgzq4ApJkwTRqQM
VBFsixLYh2WHxWyhSqoQQ6THZL4OGnj2emdHss8NHCLb9mVCyX6YOPucAu5kGysnLMX0D9Mp4Wb2ZGI3yRiJ3oxLBfQTrASXbWueBcmb4PAa//rs0DUYqzgIWeK09g5o
ia9fmNFgGjI/5LT99C91GqkjX2rCvJPaeliDag2SBkVued75yJMlPYATqw/hR2yW3dghmcK1x9mAo5MAj5zqzEVWYGeElHmQyIv6Jf/sZMEVdhHqbZnppnRnAP6kv77c
k+xUP+j7FAHOojBCerLIHH1IKEo2SdJnyzr0362qFc6onIgU92zePhfLIkRKAayqBoytnJAlkhAUaJHvWi/jRhSNyUk5VeZ7+SqbWWfc3KKAXbtaWIS3elSY6NpdD7Pb
W4t+El3yqAzVo6Ueev9Q7nGI4WDvNxZCpLNPcEFGCXQdnIYqEyr4Ne10fKBpEa5kbhbClLUIYVCxxaz3eDKS/t33cmDSk9SKNleh+t8ICqGSyv7mlCuiNFcSWG5SSuJg
h4Q0cEGG9OMNppWr1cKxYTXimVudTBYk0HRFHBbxAJjKiCbRJr2HgYyrX3ljAm2InkPELMSQBI3KYVRngPExRulocs5c9jmpgJ6dxbidcXFcgDog3tor3qUWo8jtdp5m
QsdjCaTmfg/wrR+cdLwJGeEHiLtEU2nuhPtfSEjFlAvulJ1ALzbnvAfPHHZ74+t7sVKQRByGDQIIrBrQWW+c6jZlloNdhddpYOAaTVdVPMeAH2qx/B5L2yWvUt7x/JZa
VOOFz+y20NKqTPkqx9gleMHasrD7g/DN+k3AP20kBcFDLf1xBEmw2fsUr3K5S/912s+TuB+DYKE8uJK5v+l49MqIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17
UJDn9h522Q4n5otk1oHXoSHiIPGGXZ0wMXj8mh67v80FWi2UFD4+BsyZiBKaX9JKBnkxBO53MK2SokpcypnMH43WUseYTOJjnm586pqEQkywOgRwIUYpakNvyuzq/6yr
cgcuqXz8VKFxDjVJUfNjdsyWsDqQAoaZqVJmt7qbIAeQieSRPmDxdNsR9S2zblAq8nNc4j+UG9+4Kq2Yu+vGq+Wja0Jpd8UeIghUlIpSXBGhby7SIoZ4UN1hiqBTAHR4
VE8UNg3NkkHs5eb0lm1z9tMhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbg10+KIXsFYTOG6b0aut2at7J7D5gopf3ltziTucnB4wqLpH7MUNUMCsH5HnQ2UcPZ
aa7QZ84M1Xfo1b58b77WDFxvx6iadwKbt944LUMspXFPQB1KjT4ijF3ek5qmB5wxeZeLRwEE3MinVTuLvmGoIKFJO0DeYoPlDiZS9Yorsq1P3m57oE5EP71wxv+g+4Ha
UMdul97V65UXqWOwmzgR4iPSpypZLlx+26lfb61KXBujNJIoOz+Aev97MTdhoBLZYQTc7V0V1aYBHon/5KzZ0aS2207LiBR4896tynUCIBxNrOe0POlmnvEHzG3DuAc+
yogm0Sa9h4GMq195YwJtiC7UEwkjnGxYq+DD7vjTLkbKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYiqBo+TDdha2w0Bhh+sXXRL
N3OcLkli9FN31vnndyclVsqIJtEmvYeBjKtfeWMCbYgvo5g1ut9YK0/xC2mk5Wm/LmKRiI2lIu7X97POMWrj68qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
8S7ex6qJu9C7EQjXouQOHjzwbhgEMQrcItbrsUahDTyR5WHBuhVRE8+kEqUTKhn7dkZeshZRUO4a9E3qHwVeuUmV3UcDeLGhA/7PNcP63UxB7QU5VqbUaaa46FS7cFWH
0yGRnPZE1s62DA8g752IHD9sx0H4sCfkNv7Hmh5HsnG3Pj/BKkaN6mn3eUFljDaUpkGvRgcX5euWZ+B7TtDUalMRuDicrR0NCiIO+HvoBKEJ4SnPukKbu7xhbKvbTY1C
0M9jzUA5me9lxC0sPVQPMUmV3UcDeLGhA/7PNcP63Uw+9R059eJvNX0MvzyG0DZE0yGRnPZE1s62DA8g752IHDkBOskn/alh5LtaIXu29FHP45sqZ4YalKRdnWUMnbqa
g7/lw4e3tjxkHreCiucDFgP81xEf/yCOtXCmcu1t9K6rkQl47mls1tcZmDuA3oR8GnVxUcS+eUtXy/uOTP/EOZFhnvcvzeWOvXLnahELY47kBF595Azl1vCEHg4xdyVU
yogm0Sa9h4GMq195YwJtiOP+ZSE7XaW8Bc4ewFzJBYTKiCbRJr2HgYyrX3ljAm2Id+FUBXZ3L3OKxqh0id+YDDrH/VeTr9PiZcfdKpq/A76CymdKNs4MPDwvtFZYfXzu
ruknPmnHmsLuLRZMsb55fvXgIbG2KXL7lT6fOiJjyKo3cU0ywocpNKp4zXtVHQZKyogm0Sa9h4GMq195YwJtiF+GsgSM09fsIZS7Oh0ScLEaKCOvjx0EoI3An4Z9j1m6
OSD3RRTiMWmcUg32dpP+7EwAmsMeYpW4YWfGoZsD/WlrKflcEmhVlFsA0QyL40p8meVsQA5lAgMldXYD96067vXgIbG2KXL7lT6fOiJjyKoE8rqAxlYHU9sOmJOxkfII
yogm0Sa9h4GMq195YwJtiLNICF5oJBhrWgKsWAyaM/jKiCbRJr2HgYyrX3ljAm2Il3m9A6eNrituh3tAHpYl4iraSYWNvAZcAcq4VqwxQL3bYMB/ysQAZjSpiBhUIxhZ
AAZvMxSyVxBDARl/YMiqUMqIJtEmvYeBjKtfeWMCbYgFCv0loThwzCRwybQ/hZFDT0AdSo0+Ioxd3pOapgecMZAIRH12ZVWf98urrTfYzIkA+eEqQzCWp8uMqx3XOYAK
KhIZTZze27DwDBIF7qar3MqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L7eRmbZnmhLUMss0XHltOUMqIJtEmvYeBjKtfeWMCbYicLrtqDMpk8BcgPhi4gNWR
aLM3fZDjZtLS/BNQ/WyCsAby2vpc1iIU3eKsbG/msDUGgyIc/DkbJJinnUgBuzjB7JukIBvhL6aNiYGSTNKtvE2s57Q86Wae8QfMbcO4Bz4psBaa+693yKVXWJwNX13L
SrPcvLPYyFjjYiFT9IiUB0GXpZXyFfkhDGEWD774oi9OABMmReH8C+AeZ15Vnpp7VuvRkiHiz93n7/oV2p2wsQkkCmxBas8D12jDHr5IcjrKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYgXFN8BMRtJSVeyANBcBTT0Ak/eWaZMQMNlPZIMDV+y2chHcrQ4znjc5/6r97FX5OqwAHQEw2KuVTmV0Fv1Pqs+
ZBW6B8WbMtfByuI0e1tCQOG9US/C0HqWbdazaDEyHIueQ8QsxJAEjcphVGeA8TFGbc7FMl9qAgSTTpnPjGbFZcqIJtEmvYeBjKtfeWMCbYgpoGFcLnR7LM5GtXkb10YE
yogm0Sa9h4GMq195YwJtiDpnAWVVHivKDTBw8yw4csFpL5KcJexzrz2RNIP0AFoTtCz6kGMp5+sMRbt9URKnRce8gDE803jfaXWhJiGK88ehjhkW0xZR4jr1EKYyTILN
ELLu92LMd6h28f9Lmpc9wcqIJtEmvYeBjKtfeWMCbYguX2fahGSlnU6mxCRGwGfMyogm0Sa9h4GMq195YwJtiM0IMHlIf7x/msBKJ2C747OAo79L2BhBoQd4X80WK8R1
5CJxF58DwuP+KzXN5XTAwzdznC5JYvRTd9b553cnJVayE+El44KvDTcCPQQq3uEOIEU+Did9ZGHsLn38ptmKrDenjKac2ZyKGLtbyTX9p5BMrNY5BVY5OizAUaDgeRgr
jvl0JpY8S+qpVSVJPoL7TYTIWzPbNGKz92hyIJqibP0D/NcRH/8gjrVwpnLtbfSuKbAWmvuvd8ilV1icDV9dy+3kZm2Z5oS1DLLNFx5bTlDKiCbRJr2HgYyrX3ljAm2I
d3Y0qE2B4IrjlV8NUlHbaK9NJe/7N3zFEVXzhnoM3q0ucvAcwd/tTk02wi/BWpGngg99GqT/FlQ5o8i4utgvUIThvTa4Mx1ujKr+byan55OUwE2X1ypEG6Z6I5IwXGhP
oFN7gHeT+ZseMhR+qjrtIoFnzr/WoRymbkMJlikvBBG+Rgtf+aIwriJGmjgpJ6RXcIQF6AA99K3lTtB/FTgzU8qIJtEmvYeBjKtfeWMCbYgpkNVxUjZaeTCZkezZX9CI
5uUAKwJsIJHpti3fS7BuLjIVIriuN7BePG6q9GJl5zEABm8zFLJXEEMBGX9gyKpQyogm0Sa9h4GMq195YwJtiFbi+ESrpm9S5AvBr2Su6aDeBEehDRu5tBQw9W4ARUw6
ev8KQYWvzOKCmWC5X4RSccJs2YXQA9oc7R3njFZdwbodD10Yob5BfB9SO/AapqpZgoaMIl7FUw3yc5G8BjXegKBTe4B3k/mbHjIUfqo67SI7q3S3MR2Af5WRTrnl9x/F
yogm0Sa9h4GMq195YwJtiHRwlq2Ome+MmdJj8ytzeEO34FxOCC0W7nJscbAGK64XaAneEQlA4p52Cckh9TZuS+QcCea9HYTVuheqP4K3WWkBJOmnDqjiIy9OxAxuSiip
d5Xvuzl4den6Rn/gvVwk1fXgIbG2KXL7lT6fOiJjyKoFXsElmqzjiLnUZfff/cxmvkYLX/miMK4iRpo4KSekVyIPg9hLDWvEl2H4KcARKIgnP8w4VPJT8AuTH5BHu2c6
IB0W0oco8jICNwLdxen2qwgk/t9lnCjDvmBCqlPn9AbBC6bLvtNIOdN/L+99kfCXygtO0dedXgH6lvV0yDE/UaBqm6x0xQzFXWxztp9bVfFrHFUUG7jUqde3iFySOQtP
OQkF0lFPz+ebA9jXloCzvk1/dFQI+bNoTdA3CtXKYvTKiCbRJr2HgYyrX3ljAm2IdEMpVk0/iVLB/Xc8gKO+A7ZgZQg8CPdhRMZFQ5SpNNLKiCbRJr2HgYyrX3ljAm2I
VH705XO/+qbgJyEaEzKQT2IGN0IkfcrL2dNTaCW8950y4cZoWKoLRVrjQc52GLJLia9fmNFgGjI/5LT99C91GqLp07smbLh19MGgrMxl+r5AjfzQ912b2gfKY11S1q4D
1eImKdYv44zt8lxQrS8O7iG8E+/izOgDZtCcT6SY28TKiCbRJr2HgYyrX3ljAm2InkPELMSQBI3KYVRngPExRgJM1CofmSO+4XOh3h+rI4WApjcc4q02He313LOLF1SE
beLZi654r/YQkYbBOWaLx0INjqSk8+jzkcHX3yn5PVU9bO7VZXP3hxhO7ddihD4VcgcuqXz8VKFxDjVJUfNjdkT0lZagVCqYs/29yaA+ICCKq59VLpM5SEI2mM4luCdO
azbh+vetVpT1dyPV3w1H8NE6KAgWWJvQHj1C4vHck/RQFOGxCOZLS6v5cdTMxnmT3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/ysuwInihtl4Yw6afP7tpTX
3y6FcfW3DO9iXtQUQx77Vf+2nJanp6etjaOWJJdel6H31qy+VPwjRFqTJ6z2aHYxyogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh3NLVrjjTimRkzz3aUR8npK
yogm0Sa9h4GMq195YwJtiA4w9oiG6Tj+1ilN67zao5Yp+he+VZe0K2Q2VvnxN940TX90VAj5s2hN0DcK1cpi9EDJqrCQCDOrgCkmTBNGpAwFzRp2dVdn9X0C3a46Gl05
MuHGaFiqC0Va40HOdhiyS0xz/wspaMWwXVLyrLChyXVcgDog3tor3qUWo8jtdp5myogm0Sa9h4GMq195YwJtiKBTe4B3k/mbHjIUfqo67SI79iP4oaTw163hzO46ucsb
VJ2A2BvfR4xp9dBchA0gXPX16zCf0cse3Uw7V/oy/e+4/b8P9Fa0yK+12uRSizzuVOOFz+y20NKqTPkqx9gleINxF05+fMMIhjTy+zEu7Xt8LghHoBcuEsaLLetV4gl0
5KVXc/wpOyelg6wbFq39dpH4I0x4XPfopa+G0mRPXj3P9JBE5tspAe49mi9ws8T6ujKq7Lb5ixh5cG+KtsY2C6HovsZZR/4ud/IruAjfaHU8EyhID5H/ht56af8vWeqF
WRhpwnwvXxHxhgksHVwknxbCXwVJwLPj6GenLwyySzqUieoDlwMAzd28j/D6ENZYvxe0j5Y9NEHxBvb8pP6dPvNcU1RGB/yOhfm8ZosvZsUSRqiVp9bf6hq6IpjBQBhW
4ntYDpsvEACWxr2lyAWLEUmV3UcDeLGhA/7PNcP63UwlCFo454QpjdSjyBKRU7TKB6UpWn2BrXn6MWl6FvG+vvusgKnLq+tC4WmAIYNPdvWqXU0HtT+eMVTl9oJBjZfX
c6yfIJKWjE2CEUz07/P1IbFSkEQchg0CCKwa0FlvnOrqFRnx2cZ8/vPi6/cBrmDfKH12U50T7dc7R5r/IL0e4HI73gMzvv+1OfGMEuyVGheBGsicGBkPX0c32PkFnOej
8/S85h0S2ItuLSzJw3Dng9cnimzwEO0GEmyJ6R+6ZJKNsz2djTt5Spaq1mdbUwKIh+LfsITM93YbqdOX5PjDGmHeMy3Y8Gl4gbKCmHFZPnI2ZZaDXYXXaWDgGk1XVTzH
LTgM3ZNxbtEk3Lwg3a9e1HwBsaKbAXC+3OGiD5pfLhr5Wp0NIOLUzkWuy7ht+7u0HvwXsbFdJGAcVA9TXeoOKMftUbZdDer3ETpwSK27yz6Ub6+1eb4ttUuJnFpPMlmi
kjcNPXBp4PFAtM7mq3J81ZgP9Z1TR9ASm2PyzxXsHLTrsF4E/yfoCCsMw9QlXpwfd/dbpVh75EdeTl41+3+aL0ohNJtNgnDVEe/C9LawVUQH8jFY5RCLyXnLwMtO2TuF
bhPCaJgHQmhd4PWX/OFIGWTJpIwpxkycGRJsy7JdEuZpQNc3dtROGWuWIq5SeCHZmHe529OTjppeeWYxjDul6cXWUY6udJaHG40TmQ6SxiLBJ8xc8qlPKWB6fn7Vuijq
FdJkT329i7COnhM1KYxKoYxUCyKqdgWxzULDES19Xej7rICpy6vrQuFpgCGDT3b1LNHBMbTXIInIYOl9SbMwlAgjxITbRCQt7gZIrHPM2j9TGhB5bJ0LEMimVRSC1BKv
KbAWmvuvd8ilV1icDV9dyziYxCdaU8jZfm7jVoXZJX5w70Un1Q9IUc6G91GseXXAk9uGJq+545gBhHxEfabWeP4NkIXBbYIZ0ir7hJMiMSICeZlAhPUv6FgP1FwivFOX
oY4ZFtMWUeI69RCmMkyCzcG9g9b0fPY80Qd4jJ9kbR1OQq9p3Jhj392ckNwd2iWJlPBVNowYfRoL6SVo6vdjaKcYuDT8/BCm8lRd3wQtd1wwjxEjG2g/jVWiWEFoRrQk
cgcuqXz8VKFxDjVJUfNjdsyWsDqQAoaZqVJmt7qbIAfHONJMX/pWZ9+GztYKVlE7CvLCF511yyEJHUdfjHICioCtrRvQiix+8+hfsyuorTrsBs/t4TSUAa38rHbhtiLr
lbJmdhGHhgRK2TMTZXti7dwPx0FAGBxmMHPXripzH/z+8jAyvd+6sBabQTFouHkf6Kqo9nfCnOl1hS2M6ckOJyieTFzdAmQ27upCH6zYNiItitcx1cK5ylDbiQ1hFJZG
Gv/67NA1GKs4CFnitPYOaIj0aVSxDLDVExiGWzRh8mqNcAy7OPYaHodyRIiXFxXX/Cc+TvC8YpAVrUqSFvFssj/cdFMfhkZEAMQpXAA8hHTd93Jg0pPUijZXofrfCAqh
D0aW5ArJPqq4Q3ic8Byhoq4s76+Tkz0WkmsSkzlyr/Errd+7B7GBogm4HO8GIJgk3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/ycx9wCVAdCZgFMK5RqTvWT
QNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDfvo0+10cUMbokuNWvWK1k43h1SeK32/HOTuX8dhAVQ6UDJqrCQCDOrgCkmTBNGpAzUZ9SUD3EWYoRqfNxZYsdt
SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/46Zf0DxztdDNhJSiFwGfdDoNxF05+fMMIhjTy+zEu7XuGz4cQYvd9nZbLupgYYLRH
he8Szp7LoXGyEWO45vKHIj4hCguqiTViQ+TmdiVlEEBkQqy2K9YjZeCH1DEP2Kr+xuA2z9zhzgB/7VSuVclFDMqIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mF
sb/kWnu4Yztq4q/g9gtMaeQicRefA8Lj/is1zeV0wMNPv2Nlxt/3s8GWyhfh5zyx2mLJjuGxhTZoLjjW68bX7DHrS93NrNNaX0CWkuOi53qBGsicGBkPX0c32PkFnOej
6OiZphYEvVTM/M2bKQqxrqJ3SiBZNStaEB5FbOxR1/QhjBmhBvustMO/OKf/tmILokiZvM70sM1kay/8QwD8u7nCIlu0g8zWgoHX+IvUaXLTIZGc9kTWzrYMDyDvnYgc
80s1u2OqHYTm0Fd/2Mp/6GzjyBGmNRIwfCWMsZ5KcNGEyFsz2zRis/dociCaomz94AgNDv3zl0QV75nL2CAdEfis6KSzLTlVwZ1qqThRkKHYlKH5QpEow+woh2/lKSwm
dEMpVk0/iVLB/Xc8gKO+AzYH1+34qqrVDEZC2Q4+obbw7haRU2FIPEVTdfREZzeL5yIM9OdllrMKvacu7WJvC7w0GyVjq6iKYKfCB1NViswRqLQhyN1uhVIRyPITULae
nkPELMSQBI3KYVRngPExRj/cdFMfhkZEAMQpXAA8hHShRN5eD/jWMYqNgp2QEHouD0aW5ArJPqq4Q3ic8Byhoq4s76+Tkz0WkmsSkzlyr/GTwCUN3ZL1tOOP+KsJG4Lo
3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/y7kbc71w+KajetbVReqN1RQNuG1YF0DMQaoPi6gbKncmRcNwQ7ub5FuxILF2M1GMpzploxIe3yuj9eZkQxOT6S
vCJzVEi7fQU1hJqY0xGJR/a7MB+UZd1JHic/n+t60+/tx+B7hL4We6zxndKWymIDSZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4
aqmEdkU/KN4yM0tNVEpea4NxF05+fMMIhjTy+zEu7XuGz4cQYvd9nZbLupgYYLRHcdJk9nkOFyfLPO0XPd7g6T4hCguqiTViQ+TmdiVlEEBkQqy2K9YjZeCH1DEP2Kr+
+1vWriVRPBV1Jz6N7Lw2q1TGlDJ3QcBfpMDJLF74XkZtzH0Dd64lp9Q9mHuXW9mFHx4C/O1rDopavEnM150x1eQicRefA8Lj/is1zeV0wMNPv2Nlxt/3s8GWyhfh5zyx
vg7fxSD/tPHb3jkmlyVQxFMaEHlsnQsQyKZVFILUEq+BGsicGBkPX0c32PkFnOejNEwhUCT6L9nRyOoIhVs6xTLhxmhYqgtFWuNBznYYskshjBmhBvustMO/OKf/tmIL
ACOGaEAQUR7cfpRjeJtDLS88NyVfOgL1mGSis2QW74jTIZGc9kTWzrYMDyDvnYgc/Q3CNWg9Cly6qTkokiDXWNuFhtIemJZrb2blTtbdIaKEyFsz2zRis/dociCaomz9
4AgNDv3zl0QV75nL2CAdEezYEYdoIhPdG4K27OFQYb5jiyjfzVTPXrFbZ99I+uLJdEMpVk0/iVLB/Xc8gKO+A0u14nJVQQS+qeOxX3V2Iqbw7haRU2FIPEVTdfREZzeL
5yIM9OdllrMKvacu7WJvC8Cd3b84K5sCXKusIxcsYqoDkGSLe8kPx8VxMZfCNN+SnkPELMSQBI3KYVRngPExRmNpydO8kad+8hp3O7g09RhBJmlIU7ajV4C6nYrYNjCX
D0aW5ArJPqq4Q3ic8Byhoq4s76+Tkz0WkmsSkzlyr/FZZPz3AcWNart6Rd4WnHpe3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/zkw9NfpWcXNeWQFUN7cHqE
QNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDfvo0+10cUMbokuNWvWK1k4jl3pwbUDGGMw4oTtkYtdk0DJqrCQCDOrgCkmTBNGpAyCk1Jfm0+j1gVtYW9kjpdN
SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4pXyg1SCfayX3lv4qyEiCtINxF05+fMMIhjTy+zEu7XuvkJMX5SHyeUUljVYRDEA6
Yw6USLaMdetiVxRBYN9GlT4hCguqiTViQ+TmdiVlEED+Zc02FC42LFlOtD4REgjlEvI5Z3CabuaA44eST2P6hw79tZajyFDom5bCP7KfyXISRqiVp9bf6hq6IpjBQBhW
mplRA6w72l5V0o34qZTmcN33OijE2mgl2sbCBbBI5yAEz7OH7NQB8S0bGD5jOdV7qfefUfdWnFSGoL7piGzzI/CD5FNglprGT3JDJgCOeRv+RPWUJgbFO3KTq2cRDxDh
fWFrudg4mlYE9r/LqhDYI1MaEHlsnQsQyKZVFILUEq8hjBmhBvustMO/OKf/tmILokiZvM70sM1kay/8QwD8u6LNWlfW/R8nS8UlTcov/XnTIZGc9kTWzrYMDyDvnYgc
80s1u2OqHYTm0Fd/2Mp/6Fw9sfeZjalSEPIi1hfaeCWEyFsz2zRis/dociCaomz9NYD2L1AJs9TkHn0PmW9EDx+GpYR8ADrOY6tKpzL+3RCdmay6ovqVCrZGH5f9b5v1
FdJkT329i7COnhM1KYxKoarBXwoBJykGFLECJDHL7zXw7haRU2FIPEVTdfREZzeL5yIM9OdllrMKvacu7WJvCwaG2BEPjYdOhFjTn0sB4mMR4LuQ+awoxBkqwC6aiWL3
nkPELMSQBI3KYVRngPExRoJ+0W8Uas1VwLilxtLWcKz7rICpy6vrQuFpgCGDT3b1D0aW5ArJPqq4Q3ic8Byhoq4s76+Tkz0WkmsSkzlyr/E3JmHscFqxko7reAyEluZS
3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/yAv4rZzWaJxIw+cBw45fQiQNuG1YF0DMQaoPi6gbKncmRcNwQ7ub5FuxILF2M1GMqONZCWqXKRuNdukb22XoYl
5atftZFuWsqdjA25mnqrhPa7MB+UZd1JHic/n+t60+/le49DL6G98aJyYXQe5MqhSZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4
61YI4RNJhdyCUZDoM9Ms14NxF05+fMMIhjTy+zEu7XuGz4cQYvd9nZbLupgYYLRHmy0fjgfpUFCtS7PkO0j2xj4hCguqiTViQ+TmdiVlEEBkQqy2K9YjZeCH1DEP2Kr+
COga1Gq+V9LS/y/D3AH4t1TGlDJ3QcBfpMDJLF74XkZtzH0Dd64lp9Q9mHuXW9mFP2X8e5wHH14yy9RsCd1cQOQicRefA8Lj/is1zeV0wMNPv2Nlxt/3s8GWyhfh5zyx
WlRsxP7Ej4NoqymhqFccn+xYXdrU+8vRaTlh0RWV9UWBGsicGBkPX0c32PkFnOejyYZZOJp48PYNvVe6OKg8v8wQ6sMUZJPoM6+b60gYpIkhjBmhBvustMO/OKf/tmIL
okiZvM70sM1kay/8QwD8u7O/ldGXBIvzMVW4kZd7oObTIZGc9kTWzrYMDyDvnYgc80s1u2OqHYTm0Fd/2Mp/6GdgatqFJXaJFmIkDfidZx+EyFsz2zRis/dociCaomz9
4AgNDv3zl0QV75nL2CAdEZv9AQZqT8mM6wq/ebvugE13joYKtcc7x4wCUefzRzocdEMpVk0/iVLB/Xc8gKO+AzmiTWLYHyVDA7tCIAZdL4zw7haRU2FIPEVTdfREZzeL
5yIM9OdllrMKvacu7WJvCwaG2BEPjYdOhFjTn0sB4mNtN9lD9PTBgWw5KRRSNxbgnkPELMSQBI3KYVRngPExRoJ+0W8Uas1VwLilxtLWcKz0ZxpRlIV8S4kgyxFv8hn/
D0aW5ArJPqq4Q3ic8Byhoq4s76+Tkz0WkmsSkzlyr/F6Vvdo1vZOrRVckOSW6yAJ3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/wjrI9FM7ztkukC08rcnFH0
QNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDfvo0+10cUMbokuNWvWK1k4Ie8jNRWdCPlCXS/DQqSCHUDJqrCQCDOrgCkmTBNGpAxQuxrj8/lZp/iVWaiHCRc5
SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1ujIroY6L7Q5/6ia6AKap/4nZmsuqL6lQq2Rh+X/W+b9YNxF05+fMMIhjTy+zEu7XuI2yGewAgHRVNkLO+0IEC4
8FpnaOU8oOxbgtDgG8ilOz4hCguqiTViQ+TmdiVlEED+Zc02FC42LFlOtD4REgjlN7f0zMeYYkoKnDDSR7wtQqceo6BTnm5cNYI3Vh2JxuwSRqiVp9bf6hq6IpjBQBhW
aCNty+HKZcarcFNCAp3BZOQicRefA8Lj/is1zeV0wMMEz7OH7NQB8S0bGD5jOdV7qfefUfdWnFSGoL7piGzzI9NREgBaKAQquGhPDLnenCl9SChKNknSZ8s69N+tqhXO
kXa4oqtVvNYZRPn33wM5qMK6z9P2mIN5oMzY5t8IlwkhjBmhBvustMO/OKf/tmILACOGaEAQUR7cfpRjeJtDLUIQP+5eMbdMe0dqrxkNYLjoYZX65StPHIV97J2Z3qTb
/Q3CNWg9Cly6qTkokiDXWMPxfrViDK+RuwGH77GL6bCEyFsz2zRis/dociCaomz9NYD2L1AJs9TkHn0PmW9EDze6swLJHidQq6nZT8oE1TzXJ4ps8BDtBhJsiekfumSS
FdJkT329i7COnhM1KYxKoQgqi+zc/CJS/C4NBFxG9vDw7haRU2FIPEVTdfREZzeL5yIM9OdllrMKvacu7WJvC5TQ/eJbwteIF7uZXirz2zLQDGu/1J/Ec0GOBqWrwxxW
oY4ZFtMWUeI69RCmMkyCzfu/eVKWNcYmBrgRFUSyqi5w70Un1Q9IUc6G91GseXXAZrzyjzvzqdFoZpfiV7k1lsop15xYLHxI17sD7lWXpvTKiCbRJr2HgYyrX3ljAm2I
3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/y6F3Z8kUiOzG+NIrf7hWHzQNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDdhgL4vnwr6AC78GU45bmgx
8lf0Lmgx7yCh3tMPvIOvL0DJqrCQCDOrgCkmTBNGpAwm5aqw1W+Tq18cdAINNCkXSZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLn
s8tnorsaRTNWlvawGeyKV/vibdFSSzkHcW8e+ZkZD5B+l20od+UaDo0ko4eGEnF/sjSYWEtOgAu2PZVhSK96FD4hCguqiTViQ+TmdiVlEED+Zc02FC42LFlOtD4REgjl
4Eh9vjzLAuQSLKNhK0SUP1ZT6Txt2brJMjL8eetioQcSRqiVp9bf6hq6IpjBQBhWf9tbTRCuRuc8IVkmXR9v6eQicRefA8Lj/is1zeV0wMMEz7OH7NQB8S0bGD5jOdV7
qfefUfdWnFSGoL7piGzzI011khlobcQqaagIP9pjFU19SChKNknSZ8s69N+tqhXOKl3c/Y/O2kscecbvqbIPQJ6baVfWFnCoM0S94XgfnyEhjBmhBvustMO/OKf/tmIL
ACOGaEAQUR7cfpRjeJtDLUGsMBHfMsT6V/vUsYg7ZOqXZalKGz6LvbKaQmehekmqkjcNPXBp4PFAtM7mq3J81bT56Es9m4ebg0VXf+fiydqEyFsz2zRis/dociCaomz9
NYD2L1AJs9TkHn0PmW9ED6MyQzVrVPiapWwklVHAO3gdGpV1gvEWkeFaYpKS5XupFdJkT329i7COnhM1KYxKoSyU38Qu1yg/s0ZyPN/VIT/w7haRU2FIPEVTdfREZzeL
5yIM9OdllrMKvacu7WJvC5TQ/eJbwteIF7uZXirz2zIbODdamoJqUuxN3ufwVJF+oY4ZFtMWUeI69RCmMkyCzfu/eVKWNcYmBrgRFUSyqi6/O2LnepgRGBcVzg/VXSAl
D0aW5ArJPqq4Q3ic8ByhosCfHLzfRBpE645SqfaHtKkvlW7m4NmrEngfLwII3mEI00cVAlBQIvOs3Ldb77ayrytPQgGgvhnT6E6HCAMb+XgTIHH0F5sQKIXVmyr0bY76
QNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDdhgL4vnwr6AC78GU45bmgxs94HvE03q1XQ6Do4pDkLT0DJqrCQCDOrgCkmTBNGpAz9xpNu4PFxaHJiBIQNq7K6
SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLnB0qKTRVFBkVasZ4rfLaTS43ckBNAOZ9gLIsLQM4uvk1gJM5/BmFCV37mY4767vPI
2nwprEjEJ/BEkk9longSKT4hCguqiTViQ+TmdiVlEED+Zc02FC42LFlOtD4REgjlv7ttz6sxFXvadL+yMkOh0Itga29j9WzWHanK0tEH3sQSRqiVp9bf6hq6IpjBQBhW
p5tepIjfqeJwybD+z3gb/eQicRefA8Lj/is1zeV0wMMEz7OH7NQB8S0bGD5jOdV7q91ftsTnneyk0w9Qe+3D+DLhxmhYqgtFWuNBznYYskuBGsicGBkPX0c32PkFnOej
J+bsw0iNXHBcIPYE+BwRAlKEj3lP0+QGvBwV12llX1ghjBmhBvustMO/OKf/tmILACOGaEAQUR7cfpRjeJtDLWsamCGODeAM9iMrt3+ioo/KCd0qii5hS97u1sLt5I67
kjcNPXBp4PFAtM7mq3J81UP5B3TS//BLqoDN5t8MOlmEyFsz2zRis/dociCaomz9NYD2L1AJs9TkHn0PmW9ED5ZqGn4tTX8IK+BOB91nuV8F8KU4yNrVNYyj37rNjfUF
FdJkT329i7COnhM1KYxKoc+9Y2hLuuIr6wuo4VBhlGbw7haRU2FIPEVTdfREZzeL5yIM9OdllrMKvacu7WJvC5TQ/eJbwteIF7uZXirz2zImiXnvxWEdL7GMO2TZ4ql6
oY4ZFtMWUeI69RCmMkyCzV5kFyKfSgddDR+TlMdLUSGLYGtvY/Vs1h2pytLRB97ED0aW5ArJPqq4Q3ic8ByhosWLmIJFAjV9f1zyAzuGJEYtim++Bz4208UmDu+v0Dtk
3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/y/bTKKysCecnAoyMcfar75QNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDdhgL4vnwr6AC78GU45bmgx
SPULXBh8Mkn8TAZQqLLdLEDJqrCQCDOrgCkmTBNGpAy8j1V6wnWRN1RCwqQxLnC5bj2iK1Ds8eSRrYopgplH/VOm4Dtoc6VTO9IgwMUbG1u3YfZ+V+LRwUs10qucagZo
M5GvdOdtdaoxjV8jnJBiSoNxF05+fMMIhjTy+zEu7XvaVRIf1dMRFCyqGnRWbzgi1pUT1gtruzDL477SIj7rWD4hCguqiTViQ+TmdiVlEEBtHSTLpes4HhzMSie4S5GK
zv3QzTAeIyxnXbAs9MR7XuPwSLf1NzWgqmvdjD16+hltzH0Dd64lp9Q9mHuXW9mFVkvdnPlMV+hPEvHP2TDFYuQicRefA8Lj/is1zeV0wMMEz7OH7NQB8S0bGD5jOdV7
qfefUfdWnFSGoL7piGzzI2b0RqDJT+CEUGPK86mBSU19SChKNknSZ8s69N+tqhXO5yiigsWAFQDeBRfyPBO2pbFSkEQchg0CCKwa0FlvnOr7wKTp8uziRn2+XlMRgYxd
KkqBG6sU/yv3GyHI7jbzHcqIJtEmvYeBjKtfeWMCbYjTIZGc9kTWzrYMDyDvnYgcuc/k+OXiweAW5ELnA4Vm4FOYpOXVZtX5padaMFZXfFeEyFsz2zRis/dociCaomz9
NYD2L1AJs9TkHn0PmW9ED6MyQzVrVPiapWwklVHAO3gLjbt3LCvhGuxpqFWxl4p/FdJkT329i7COnhM1KYxKoT65JshVNzd9hY9pNxbeZV7w7haRU2FIPEVTdfREZzeL
5yIM9OdllrMKvacu7WJvC5TQ/eJbwteIF7uZXirz2zI5ddGSy5Vebt9KjXoQ5wBIoY4ZFtMWUeI69RCmMkyCzZY/ET5fs0qnvvkrETVf2KzSgkK0Osz/h1YY8fSHvauj
D0aW5ArJPqq4Q3ic8ByhosCfHLzfRBpE645SqfaHtKm9yCBcufzOzHKFnLvMgOwTua+/cUr50fsNVaCl3J+3lytPQgGgvhnT6E6HCAMb+XhBQaZvjjr5tRtGRL1y/ASv
QNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDdhgL4vnwr6AC78GU45bmgxOHvturvS9SNunUDayby0yUDJqrCQCDOrgCkmTBNGpAxzSNHmeCmpSVxpGSAsQ9Ta
SZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLnI+mbLpUpSBA0tIDiCHBRLI3ckBNAOZ9gLIsLQM4uvk1+l20od+UaDo0ko4eGEnF/
CAxs3hkbUNr/LLllFsdpnD4hCguqiTViQ+TmdiVlEED+Zc02FC42LFlOtD4REgjlB6bzFal5+y/XT5pDAUshFbuRkxvR8jmt/P/uHxXrTJUSRqiVp9bf6hq6IpjBQBhW
1KW8srTCbx98A5MV2pi2COQicRefA8Lj/is1zeV0wMMEz7OH7NQB8S0bGD5jOdV7qfefUfdWnFSGoL7piGzzI4F+WB7OU8L25ayuI/1oxuN9SChKNknSZ8s69N+tqhXO
NrLV5s7QPXFw03rRqO9XIsWv7ey4BTkHK5Ak34ofE4khjBmhBvustMO/OKf/tmILACOGaEAQUR7cfpRjeJtDLZYHDdwxrrfJbI44B9VQdVVkMx3YhgY66MD5qJ5f3b3A
kjcNPXBp4PFAtM7mq3J81a6tve0DFPWXXGGJmVLbYN2EyFsz2zRis/dociCaomz9NYD2L1AJs9TkHn0PmW9ED6MyQzVrVPiapWwklVHAO3g2UgEIysDFn9ucT1KiBklA
FdJkT329i7COnhM1KYxKoRy80jEg131zs9VnjcCI5O3w7haRU2FIPEVTdfREZzeL5yIM9OdllrMKvacu7WJvC5TQ/eJbwteIF7uZXirz2zLCQnlTjwqg+lSdQMiNIMQW
j0byxz1Ozwgny/kA+JO/jX1sQXCmnRN3dSPNOn8Ykz+LYGtvY/Vs1h2pytLRB97ED0aW5ArJPqq4Q3ic8ByhosWLmIJFAjV9f1zyAzuGJEa3SbFzeHs3nbuHYO60ghsd
3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/z6QeYg9WrK8D5PQPobWoRgQNuG1YF0DMQaoPi6gbKncsDlicVnrgUWDK9VOIDcHDdhgL4vnwr6AC78GU45bmgx
EkMpSPrruZyQFoIzqTagykDJqrCQCDOrgCkmTBNGpAz3sHYl6ELGDojTVKfNKHLYSZXdRwN4saED/s81w/rdTFOm4Dtoc6VTO9IgwMUbG1s1Vfq2SA8Qzh6XyHmrFSfp
3W0mzfqhJn+IHnJip+g2dINxF05+fMMIhjTy+zEu7XtQkOf2HnbZDifmi2TWgdehOaGB12kZmYTpt9InSB2QdT4hCguqiTViQ+TmdiVlEEBtHSTLpes4HhzMSie4S5GK
11h89KJzQowa+5pSzOOoLcqIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mF6X0dijAimjUaP5li8bJkVOQicRefA8Lj/is1zeV0wMMEz7OH7NQB8S0bGD5jOdV7
tZ2SSm/teQqlvkjh/dsCbB3xNFk3tNezh29P5W30qomBGsicGBkPX0c32PkFnOej8Dc6RxBSV0Ag0skXdMphby5ikYiNpSLu1/ezzjFq4+shjBmhBvustMO/OKf/tmIL
wE5wpFI2s9yjVgXmnA/BX8PxfrViDK+RuwGH77GL6bDTIZGc9kTWzrYMDyDvnYgc7CAGTtCECKXBBMEApE5Us02s57Q86Wae8QfMbcO4Bz6lEGXn5EpV9CcofEFEDkTv
CcBvhCSt5lzzPQLIGQ0EpsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IeR9uAooWsrumTiNUSxyQe/qCP+E9anMlIyBnau+rmnXw7haRU2FIPEVTdfREZzeL
/uilzDtVzG/v2wYdM0SdBcqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IshPhJeOCrw03Aj0EKt7hDi9HNo0x8pyon7YRDuq2GW2ZcEP6LjJYOZ4ZfQlMiXDk
v3GDVd7dlPliFVCHKyNqyQmhzrVJyakqL6ccJIDeVvjafCmsSMQn8ESST2WieBIpcB0PT9BrXRqvz13urvxCHpTclEhZAeSBh0Y/zJsKWbsBX+AZzxq5GYQFvz4MUpaO
T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCAehBwnGTvkcR99Of78esbuSZXdRwN4saED/s81w/rdTC++Y0NvLvfRuoM11qesNWeENF86I5xLaJXox0D2qzdF
yogm0Sa9h4GMq195YwJtiEDJqrCQCDOrgCkmTBNGpAyPz5BBRGSTdiE58l2nVcALQSZpSFO2o1eAup2K2DYwl5gZxeMUsMkFl3JFLzm4UYFrg6qWlqhoJ+zed+WI2hpL
ugSHUx0t1kAEhXJrUNlTrXIHLql8/FShcQ41SVHzY3ZE9JWWoFQqmLP9vcmgPiAgx6ObMz/SF4CFSGAaCUQUcVyCXWM/+e5NkUlgBSS4HIUEOHAYSUZrnzoCECeKvZtG
N1qOuyQmPmCKB8+i2hMab5ewoIPnpv53yku49gQU9xZ0QylWTT+JUsH9dzyAo74D6WVftVpo0KBgc38BslIMI6felt1bZyAt371qIqTvO0K84i62FxEvwhRtWQh9Ujdl
2DOuPnbzdj6+D80OM99v1EINjqSk8+jzkcHX3yn5PVUmuuo71aMyaeAxdGIkvTzlwXs9S41M2oflb6dEEB0+moqrn1UukzlIQjaYziW4J05wKKCVtSyPyIf9OJFmxAG8
6xy8+IPZMHJ3jHZ5TerZT8qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2Ibcx9A3euJafUPZh7l1vZhbEZRch3sVC/KwHqluYdB79bpj7Hr53P/Gq0aorMZqR9
SFUpCOymwGPW7UrFoIukUIfi37CEzPd2G6nTl+T4wxqf+SWWJUsyFnlGIDK0qiq0NYa36SNm8vnXng7b66Wt4d7TLRmxdYRpn9b++ETtzI/hsgeBRaLW5blz0nv6+dao
aA5oCFAD2IqjxuNNpJxkFEibMTS3tbTrID/469ex8AtkyaSMKcZMnBkSbMuyXRLmMut7W/ytdkjWxkAxIPlzc9wPx0FAGBxmMHPXripzH/yxq811Hos2wOnqPiXb3uRt
rl6GzEjFrToJhl3WfxMF922v1fa3n2hUJWA8P5OJGLdwZHhgTEDLa/eFu7mZ/CbEKWfX4vprmOGu8srb2GbEfP2tn0rZDQHp3KRLDJ6DcNgkIqfK45Bkr7qx4YhoBfqw
3ZxRf6QF3YOhXQCMrdR0vZTwVTaMGH0aC+klaOr3Y2hxoBIDECt7ah5rfIQ9HiF7eTpWnkM9e9qRS+W2ldBabSGfi4E2fLVLy1fN9bMBs+3zSzW7Y6odhObQV3/Yyn/o
BkH2SP20kbDpu/TWbBX9gsvc963oqGA6BeMEA0oAppxt3WE729ZK+LYBKpHOlbHk9Vo12cYwFWYgikEuMEmvWsqIJtEmvYeBjKtfeWMCbYiqXU0HtT+eMVTl9oJBjZfX
XwGqd55mQiP5EUFlmC2XW7FSkEQchg0CCKwa0FlvnOpxHkbPKIS9iH9bielhvGtfB83g+X1b/20MWatO2nF7yVKTrxHtnWxBqOCkrQb60HyDcRdOfnzDCIY08vsxLu17
r3BHxdEdPsnrYsA3HT2E8L7GHktMUlHHsWDlTchce0hqomAJPclZBfWv/JSelZJ3XCaHntcoy8MWPz16fh7i0mTpf9nHsfAuhtxZXQA2aujKiCbRJr2HgYyrX3ljAm2I
HnxxE58x7qzsr23/eeD5yt4bKkCydu+bhoGAWX/VJZNcNTOtCc+GcEoyWXd2sbjuYrVu/YCaUWSjIu+r1S9bcyEZIWS6VRyStpTqCI/OYmU9byeZFLWBz5MiOduS6koF
oY4ZFtMWUeI69RCmMkyCzf4B7vWVRFfGSWCrUbdoosjkpVdz/Ck7J6WDrBsWrf12AjylOwG6aqmAiWEfMYVrWK86srOoV8Nc7iBMM6b6PeiQieSRPmDxdNsR9S2zblAq
TBgk3x1l/3O9DLMjR07PJ24TwmiYB0JoXeD1l/zhSBntLhF5lk8tVI+Enocprf5J5NFUvvQt2QMl859chhXei5d/5XoLnJ62fHG7YFQ/C0zDDkBpMMMuC3aEyxQL/uJA
ggHvRQlcOeGYbmU9fpnD431IKEo2SdJnyzr0362qFc6Ic7/FLbUYQnarhH0YPMzMDt/p2Jnotw+tvOsjV2PhPSWIRGcXkbMyDzesxELzAagx3kMlFcImKmPJ2rkD9ppw
qZHuNmvGrw2vK/JCmDmLva77s/BPK13KhyVRPG2xDhc8EyhID5H/ht56af8vWeqFR8M0Wz797RkQquWqd+oRNUmV3UcDeLGhA/7PNcP63UwvvmNDby730bqDNdanrDVn
hdGjW52EIvIfw2vdC99BIMqIJtEmvYeBjKtfeWMCbYhAyaqwkAgzq4ApJkwTRqQMQ8e4Y61PFrQPqpH/0QFk0jLhxmhYqgtFWuNBznYYskuOEeq51Jn2VxuzCmHvwpvo
aqeZ/ji6C+nvTkMaVjfCI3DvRSfVD0hRzob3Uax5dcByBy6pfPxUoXEONUlR82N2zJawOpAChpmpUma3upsgBwZEG+A2CTidlB3wvHMt/bKS9p/Zq6lLEXw1tS25nLVt
UfiDPcrHEqrsRqcRHmEteiQX12+gjaYCBNR5QcsJV0jKiCbRJr2HgYyrX3ljAm2IFdJkT329i7COnhM1KYxKoSEtpyJzxUvTubbO+dNMWvqwOgRwIUYpakNvyuzq/6yr
kgNoJd+djeZpWp2KDHasqRt+KEDPu5URuDIIaTga4FxcNTOtCc+GcEoyWXd2sbjuNmWWg12F12lg4BpNV1U8xyv7Z5piUGdNYHFs6eY1Y71TYyTerXB0su1jYcSlJ9gi
PQ2gTXk2f+JQ2IhokUeOUtlCV0UafUhRzM4chONDFDD+WNCKwabbQzJjx+iJHz5oes1KdkpWhNtbPqjqL08v+BJGqJWn1t/qGroimMFAGFbbmNjAg1IYfBpCGrbKiFQk
dKmUESfDBEenzRrN96eKk5jm9c83TV1DjxvZyJWcqmiMSwX0E6wEl21rngXJm+DwRlhR6QicpDPVNeJIOAWLYOnHVftzjYQ56eym/QM73ELoCUJ/yXPCpBCp3Xouux3f
E7rddoogtB9oG/8HLCS7p/gSBbmfAKsa4sxEa386Erq2lI06FVws7R/e0mm0UfEWKnIMB9KcfZHV+WmAiMOGQbUYQ+P0rmzZG/ob/OOlmIorT0IBoL4Z0+hOhwgDG/l4
7xNsfSnawPp0418jdqIPWAqOyhoKxJaGCt4myMNaNZIVyrvKNuQLuA5okizpZqbVSB6jnxB7C06R0m4uR2cisvNcU1RGB/yOhfm8ZosvZsWJr1+Y0WAaMj/ktP30L3Ua
qSNfasK8k9p6WINqDZIGRW553vnIkyU9gBOrD+FHbJb2h0CgGGsAmKr1gVPQ99p+zvlkrhGs3RdsCM4G6GslFCJdTb2+e5138jetHbtSKOh5lx12gS9Lt6ez+6nGw0Bt
kjcNPXBp4PFAtM7mq3J81fOP4rxMx2SMOcNT24JnUJU2hoSNU34eBz9R/XhY8hxbbd1hO9vWSvi2ASqRzpWx5Fk6ofNhz0GeBRaUDKdlD1ZP3m57oE5EP71wxv+g+4Ha
ql1NB7U/njFU5faCQY2X1xnzpDzanRKVU22bKyapPHpNf3RUCPmzaE3QNwrVymL0xARU36a2APFypw3tFicy+188mo/y0urESbppdTOxcTCLYGtvY/Vs1h2pytLRB97E
g3EXTn58wwiGNPL7MS7te1CQ5/YedtkOJ+aLZNaB16HUDpjjNeqx8Y5CT08ugsW9aqJgCT3JWQX1r/yUnpWSd1vNAhueOdBJ4tOcLDU7Zb/TeA/sB5NfWDiRKAQGnPrV
yogm0Sa9h4GMq195YwJtiB58cROfMe6s7K9t/3ng+cpAcc9qtCKbhqQ6wJcJ3tYjyogm0Sa9h4GMq195YwJtiJ2iGb5ygLoL+L0830K2QSfAZ/WU0ctmSBVnMJqR45Lf
LmKRiI2lIu7X97POMWrj655DxCzEkASNymFUZ4DxMUbpaHLOXPY5qYCencW4nXFxZEkljiuTsidH93CjhXspED4gfLIz5h0+K0oXuKhg9TR9/qeu2Y67DtcEG/yNy/zV
SEE/RIUPM/uKy+F7A5BNIWJVNCmPIBFaSqGHsvUMjxRFTtzj4ByygKnyQoSrGrIy/F7fKz9nsDQCTNzTNI5APyYAxS2Bjw60RfNGOilCBl2HovDWMMl5GXoICOelD5+T
jdZSx5hM4mOebnzqmoRCTDSXFZ5fJwtpSZ2s2O47T9mBGsicGBkPX0c32PkFnOejSHbZCEodin2y9DUr4EHWF0R5fAOqRMZI8caN1bbRFZWA3DZOzf2yZgWUVoD2GRCm
4K5PcKowuG+hZ7IufxMKaYgNGvoXOVOt4o69+hNKIyi5FYt8YrWlgrxPqP1u81KPeZeLRwEE3MinVTuLvmGoIKFJO0DeYoPlDiZS9Yorsq2jJ2f/BWdlPrqav0zEHAWS
VO7qieuy4n4oKGRUjhx6HtxNVTyrJcJJNJwB/K0ICjVWapOQ5OY7MWfmsHTheYcSGfAdtam0RKEd+xZ3RrDNhgzSynTfQGXOyzeTqkkBffRDDeD0j3FDeVGlN1qtpata
8iRjvq0o0ZdwHrs6rDRshd+xI+G0hm05bdTYTpnr8nXnIgz052WWswq9py7tYm8L4XNyYFjl4ut4c1xyQElywNchdOHU/fp+Zqxg54D48QTNESxCKa3fkie2WGzq3TkL
SW9NF6CKBuHLdrfZ8dEq9ryXXHZzsBb4uHLOBxk5GGUwfBKcUi827xExHJIK4liPzSU+SAcAXhiVU6sk91xVrsBOcKRSNrPco1YF5pwPwV9sqBMZ5IJ9uvwq6fk5JJ+T
HsgtschURjQM4IlybnR53wyEbC4nQRjazlycDJdkGHfATnCkUjaz3KNWBeacD8FfyaAg2UBSNt1KI2pwCQU0/BRDAnP3f+H43uGDCmfEKAbdKpH0i4bH8uAJY/pXzfjJ
F637nXWg/DhjAeLtTqzIAeTVDMkkcX6v4RRSAA6tC2JVAtaRdzcVQ0ua8Z7B2BO4v5ULOlt8QBoVft1iP22YZjpOeuF1Aekwg49T9LLqYTvL8iCVJIv0H6UPG/f/xagL
jhHzMmF7eRz5kBd7qcgEttZEh1sKe8G7v+ibGV8Rqm9sSNnxWto7+AzhdjpJcPLwJNhv61neDU9fOxEMY1rCqW0dJMul6zgeHMxKJ7hLkYrHUFPVUrZY2j800MxyjiV0
B6x6jnv7FtSRCbHp53CDWMAKXX63Ck7+j7kx6Xx7Kx14hHNdE0gTNC+PXxrNM3RS97xmSgVZGZOhzNt6OaoCON4mtnyJXOqU4sjfHn3pF7jACl1+twpO/o+5Mel8eysd
bDI+dBN7LTGb/5peFZZZS5GPzbOmy2Eg8tLWuNL8iPhtHSTLpes4HhzMSie4S5GKx1BT1VK2WNo/NNDMco4ldHwoAEmBwRQijdxP+k0jVwok2G/rWd4NT187EQxjWsKp
jriEUaKCbNLG/fe/9dtJlfCSi7nB8FjB06Jmd3bWyE7nIgz052WWswq9py7tYm8L4XNyYFjl4ut4c1xyQElywDcOV9nZe1ZLDVGK3ebwrfTaqSQH0rzJWmJSnR3JLNF8
htI/Vu8MJaYwqhb4WZAsFNJuCqPrUf8pcF7jSNahz7FmTX2JdZhfb35fRgszZj3S5yIM9OdllrMKvacu7WJvC6V/H4LC56YqZpLvuF/eEFeU2VIwjw6TFq9V11Zxkcu2
rDgcaeznJM+WtUtrnWcd3HP0X6OeaOViqLI7IZ78qBoYvxg0/eo5ddIgHhGP42Puv5ULOlt8QBoVft1iP22YZjpOeuF1Aekwg49T9LLqYTv4qWhOzVsRrYa1g8lN9UH8
SW9NF6CKBuHLdrfZ8dEq9m4t1W2S7Ifz0QWIHH6/N3LNJT5IBwBeGJVTqyT3XFWuwE5wpFI2s9yjVgXmnA/BX9eMDnZigfh6L3mW8a8jri/FXeSGmDWkt2iWwF/WSGNj
i/7P8e7ESyfLyrpYbp24YhVjMktaXGVBTCwoFBlbaOUYvxg0/eo5ddIgHhGP42Puv5ULOlt8QBoVft1iP22YZjpOeuF1Aekwg49T9LLqYTvYQYQnDrfDJWnVOOmFCiN0
RK6q0VoLiyzL4hM5mmYYx/oYrfj5rhAXr51xMwgVqNBbFhvDE/8zqWE7bt4FH80q3SqR9IuGx/LgCWP6V834yRet+511oPw4YwHi7U6syAH+xmWhazjOQOBOIEw0Sh+M
5yIM9OdllrMKvacu7WJvC/sb8+0DtJYJ43DHF9xz7oe4T1VUnNiA3TAoF9UK9E9I3SqR9IuGx/LgCWP6V834yRet+511oPw4YwHi7U6syAGxN+4jmp47gFHuamunQjE3
r3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWdAe/yNrlvMggIHdIJ7coJCiEUPjDsssWg1Vt5Z7RbKOEquAhTE7XoORyUg3wBK/+j/WjxPbB+zCONnzyOHdWt5
v21DjKfdvNjMXd1nCzho54bf8DVrIL/kBizjLrELUq/dG33T2WTp3w6Xufevs7+ikaUI6BdDB4cBakAqvDTW0srOfndS1iyFM5PAOFIyQpQ6mHABMu1oDkLQSgigrVX0
OK0b/Ynjx+AVPzpDcfJmm/+q5nY7WBv2SyrLHBK7AUhI1mh1FNCh8htDhUnJ/pgZsuGgY4ulq2aX2YKDLM1hI/F1qA5EOM/7gQ+GnxdjiLXsI+cQxcBggq6uR3sFl+AB
h1mVRTdQuGXbKqXcRIbxHP/Di/Ff+Z9E+2JRj3LZLxrDThk0HSbbuy/SuJkQkbxpBWg8Yv8Q+rv1Xc4mASTaftZA3k0EnrdhFInzGNbJ/NyfqJ0U1ONzIZ0WhzGMWU2y
Zmi+bIcColL92oN3iK5Iy91t7KWr0BjZAo9MS9mY4oItcng616xtREqzh2+vbdIBdcC6FGI5wABI8GggYAmeigEFWBYWc6Ue1zxHl6BbIVWBKJojEQO7BWGosI1j7H7n
NxOy8/FeTh+XXRkPlltRH31FKE5fikB3n8aah826wa/xZgJA57cczZTtM6fnsWM8rfm25nZwMmGz+uYOnQ1be1pOoFOQQhy9GXJy9yVSq5opDQdEMd6RXVsMJI/+v0pE
Z3JCNYv2zsw6O4Y3Fh11pzmSDmgE1eVmmdPvwFH0mvqjfsWuKq5lr+IihlDWJbcymlABHxVEp7qK0GFs4OAdwmdyQjWL9s7MOjuGNxYddac5kg5oBNXlZpnT78BR9Jr6
o37FriquZa/iIoZQ1iW3MkJNFd1FE48w9SeJ7UZffgoDzUj32VlmfBOUxtFvJU5wDmlC5SuGORuXNB46ezok/nVzWclE087CW6WrMnOpGN4QekTX8fdxAXvxfOqfUEVt
Sq4CFMTteg5HJSDfAEr/6P9aPE9sH7MI42fPI4d1a3m/bUOMp9282Mxd3WcLOGjnKOoMhv7QyceEK1lVb2kOW4I1nolwgOErLBgSZLetOuurpY9OqzrTG3VR9UcCk3LY
nreOuqgKTuhm8gA8sOhYIWrIrzzIZ4liGaGdfJH4hNHIeNA+qSDzS6dpcqE6TmaiHfhfdeTx9aNqPtrXXY/6/A5pQuUrhjkblzQeOns6JP51c1nJRNPOwlulqzJzqRje
IrSdQm+FrShaVenAAMyR3qtMqVUx2kbcRYnUB5dHWgSrpY9OqzrTG3VR9UcCk3LYnreOuqgKTuhm8gA8sOhYIWrIrzzIZ4liGaGdfJH4hNFtAVvoHg5H1UOTAjc5Pbi4
r3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWdAe/yNrlvMggIHdIJ7coJCpQk27gt2qyUaeM1gMTi7UrPR3uURSNWzbzcV8PIfbtrSBoqsTXZBfKS4CqWNm/17
BobYEQ+Nh06EWNOfSwHiY1JNF6P4jjkcrSioL7yu0W4ZsUXjwz/aOzuZ523TzUbaq6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCFqyK88yGeJYhmhnXyR+ITR
jRmvXzunehtEIJ0XKYlsSnQPXXucoU2GZEUGoDIlD67SBoqsTXZBfKS4CqWNm/17BobYEQ+Nh06EWNOfSwHiY1JNF6P4jjkcrSioL7yu0W4aICDJpH9pFt3w8BGphlzc
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mNSTRej+I45HK0oqC+8rtFupJ/IJMH0/EF9qjmSs3K8j7Uj3o591qmt/ATeh7mZ9NiHWZVFN1C4ZdsqpdxEhvEc
/8OL8V/5n0T7YlGPctkvGsNOGTQdJtu7L9K4mRCRvGk5nT2MoW7eoPZqELqbhBKQtpzsxfRgVAH0LvQCU/Sx12j9cy7XxalrE4vLfskOs3pAt9w3BZXKqVM8UkrHqlw5
nomHSygsfSVedoWwguqkkjFdw0l5g/c0hKSKUhxI/Hk0Yuv0O/po2woqlrVBpjasJ6XLf1I1w+wWExAco5CwZrqo4MVa0I9vRufFLah8e6yEebD0LfGTnjWLHEdIe997
h1mVRTdQuGXbKqXcRIbxHP/Di/Ff+Z9E+2JRj3LZLxrDThk0HSbbuy/SuJkQkbxp04ZaisF46KrT13mh/tmJaDFdw0l5g/c0hKSKUhxI/HkCBZ49Fb1Xv9wjvkNawxdR
+Z6bBjDSN+9fJOKVp3I8En1FKE5fikB3n8aah826wa/xZgJA57cczZTtM6fnsWM8rfm25nZwMmGz+uYOnQ1be2pAxxHkF+NcG+7tih7VJQY9MI5bQvq0DRFT9Sp/3zYu
aY3SecHz2Z+yApnqIuEE+GbpryntX7HwLHo9PhKV0X5t2V+Dl4Ws4gJo7lLSpMSTW9QMhXWvXDtU+RWN5H29YlXE0ARTae9NtROUTI9Pij8xXcNJeYP3NISkilIcSPx5
b9sP05/y3G+AHtLYUzCiz7wP4fqm5AFuo6uygV4dlWfkaDRMoeUog81+PEF/MFklkkynGI6H7x8q+qn9hnbRJ/JjfwbzI/zvDL9geEfJrdfkaDRMoeUog81+PEF/MFkl
kkynGI6H7x8q+qn9hnbRJ7RfyZdUQoi+7dOo/WBJaV8W8L9zKzQ3ZeLeMA9SnAUK3jKqZr4lPhU/bmRvaQEyRoXcz9LWnjX7aM1FXX9/lcFff6P1Wbxq09BJfnweI1uE
XxhULNHYXaoR/kCmXPnSUqgvBTfE6ZxP5FSyKZjSpCU1X1NRH9sxEmpdvhN/dvcic8zoOFdJccteiSMYYAhtBp/ntXmEZs8SNiAVj7UC6+YyvQ1z0lbgYH1o0CmLcgaL
bUBjdYThPXR3hCkBz91awG/bD9Of8txvgB7S2FMwos8EQP9aGO8GEjV3gLsobTLEQ8wYiMQYLpDIv/lkzfo9Cl9/o/VZvGrT0El+fB4jW4T4eGkqgo9aeUoFzBhxo1L+
SBhMCJ2ybDMtLcywzSeDR4BLgHFuHYVmGPlZlXZtEk2MD++Pl85CSlBz8ryXYSDlq6AOZGJvlT4ZTA7TD1Vu+YI2o/SutWbP5/rSoMxdU6fi7e5bvtLrG5zFiVbm6AVu
jQxezLAs8fWMyykcrQSAdyg+vrW9xFhmrvHetGFVZI6z0d7lEUjVs283FfDyH27aVdmgwS2YE7P6+awFzsnab+puZbMqUPQUSOtNQjVlGfc7DAadA9FLJYcK0ytMuHlN
FvC/cys0N2Xi3jAPUpwFCno6Ofr3EINyGUbjDnLoSG3aqSQH0rzJWmJSnR3JLNF8BBrFAGOYrl4uarK+eCfXgtNvRd5ZcSMacEf4weYzhOZWNhi82WE/OvQ+gdQ7O2WU
bKgTGeSCfbr8Kun5OSSfk0bwWS4nDUYA3Orym1NNB/+oLwU3xOmcT+RUsimY0qQlNV9TUR/bMRJqXb4Tf3b3IjP3Fcl5U9gLCT9ugjg5HaPt7cP/1aPSVp/7c0zL/PeP
yqI8gsKkGbSHN0zuq4NphNqpJAfSvMlaYlKdHcks0XwEGsUAY5iuXi5qsr54J9eCOq42GxPYwW0EFJZ1AonFrJ/ntXmEZs8SNiAVj7UC6+YyvQ1z0lbgYH1o0CmLcgaL
5SrV4yimL4mojk4mMvOl+aTMqoKLZfVPI4b46cmqzueWq9/sI/bKKhiTMxVfAYwb5Gg0TKHlKIPNfjxBfzBZJfRmU/p2Df8c3brEJvJLtU1IleGQ+M+RS+93y8BhuTFv
3gviT5Rm++4A+a/sW24Ll2ykesuufs5l3rjkKvHC+YhLDfgYG24JTKBgYv6D2OaFU+STxei6UL6dy+Zlm8ttkoccY/1EMLMTNlYvdE4bXcr0Uc0c0Yesv2VgY+TRMRNJ
X3+j9Vm8atPQSX58HiNbhDEQhcDcgvTvDo/hp5SqtFDwY2CTKtYtQzC9wwECag1m0XXLiFLC8esoMhW5P0ffwuRoNEyh5SiDzX48QX8wWSXvnnD1ZqPY2DmsgaWQEO1x
MV3DSXmD9zSEpIpSHEj8ebhcGHDNJTMn235+j2G2oe1IGEwInbJsMy0tzLDNJ4NHgEuAcW4dhWYY+VmVdm0STWDnTKwI90v+se7HDadd2iTbwSjFOR/izcPBStikgJC/
6cqFMhGP6kgIoJuqCGLb/W/bD9Of8txvgB7S2FMwos+4hDu+y1t2utWiPIifJr5cpMyqgotl9U8jhvjpyarO53KNwfPwGwmen/+LpcvilgiNDF7MsCzx9YzLKRytBIB3
dBxZXw74L3bLhaKWTV7gMdqpJAfSvMlaYlKdHcks0XysfO78/EDPaGj/rB02vDVdSBhMCJ2ybDMtLcywzSeDR4BLgHFuHYVmGPlZlXZtEk1QYytiHG2PlkYDpfh9kURw
1K5w+SKFUjj2U81G0NGKnCCBAu/ZH0Mm/PSSPjUPzW9v2w/Tn/Lcb4Ae0thTMKLPg4mHQ0Clwh3kM4i7Lur9k+QB0E1yDpjXeJCM4exinJOmEft8lmo2B2eECO4OItQn
VdmgwS2YE7P6+awFzsnab+puZbMqUPQUSOtNQjVlGfdzLYFpE74hg+TZIYTFc2bgEQ/T7p1kjZyHv4ZgoyCwmDo+dFA+xvRrIPs03BZ+mtEhqAeWYwN/W2i/ykYyaVcw
bLHQf7AsEGvBCTmWSwjdA37mjNwMr9U/qfU7hfYmN+0z9xXJeVPYCwk/boI4OR2j7e3D/9Wj0laf+3NMy/z3j0lNdZGroFpITK34r1uT2AqkzKqCi2X1TyOG+OnJqs7n
tKXEdLgHQuOwWj1nX7zoGuRoNEyh5SiDzX48QX8wWSWilbH7jXEw5Q+2ZAL3ADuYjjAMUdWiXWdX2PrsAmSS/3X2/dtOtJUY7NzMKaVcjjMLQER1CMLWWbziaX8lzI3o
TGWABKCVUEkIXPfXECKvh52JZrIWCisdVRIxwCDaV1jMT5J2BCiWisQhHmxYCjoHRK3bHI1IXhexJGtBd+VwQhpwjgfwAbLWGDzzFUkWxH7qz755oh5ZT7lrQb0MBq3/
IB5WfAkvbcUiQjtFnDAgF1ebx0isu/yfCvfhFVYaZy13fxX8o2BRfh4M86HnCqb19dvneaEQqp39UQ8p/B27o8kFEbPXYniJyOuQJKYbMIBwn5qr6wIAzof/KayrpiwN
V5vHSKy7/J8K9+EVVhpnLSksgHaxWJUmGGthPi8iGxZBep2UAxchaHIq4s+SnPbLV5vHSKy7/J8K9+EVVhpnLfnImcUAuaTLGT2zBuHnILlWNhi82WE/OvQ+gdQ7O2WU
Dkujz51FGLB/LVJOr3+Ok+1OHRxYRTSifXsa+Q+C5vBWNhi82WE/OvQ+gdQ7O2WU9Ijx+1keCvDu+MCJGXPhCDo+dFA+xvRrIPs03BZ+mtEB4LF7YWrbL5wdKCibliRQ
PuNMVqqjaZ59ijstJ3PQH//rs720g1p6feJGrbWpXNX9w5Gwv76d82EwCnKeOwrjXDIhnBy5TEwh8TtfDv4ZppozMh/z2lr89ERm31kdOyOO4rKyOKPjkiW6f33Rvjka
fUUoTl+KQHefxpqHzbrBr/FmAkDntxzNlO0zp+exYzznj5pQLKqgs6BhXQqQjjNxvA7BxmkPzzM26aP52n0WXjRi6/Q7+mjbCiqWtUGmNqwnpct/UjXD7BYTEByjkLBm
ZeqZ0Fnsxs0jzb1Lv5dd/4pDHbRSJfSWriYF6wz3KD3/quZ2O1gb9ksqyxwSuwFISNZodRTQofIbQ4VJyf6YGbLhoGOLpatml9mCgyzNYSMgHlZ8CS9txSJCO0WcMCAX
tpzsxfRgVAH0LvQCU/Sx12j9cy7XxalrE4vLfskOs3pAt9w3BZXKqVM8UkrHqlw5aPCCyUl+u78p64E1l9Gf1aulj06rOtMbdVH1RwKTctiet466qApO6GbyADyw6Fgh
asivPMhniWIZoZ18kfiE0dTapm73xXdR12SWxHZZoFL/quZ2O1gb9ksqyxwSuwFISNZodRTQofIbQ4VJyf6YGbLhoGOLpatml9mCgyzNYSNOiSmZQZtWuYM6bxgzLkJH
KQ0HRDHekV1bDCSP/r9KRGdyQjWL9s7MOjuGNxYddac5kg5oBNXlZpnT78BR9Jr6AIqndAjYrJ1Ji1nLFyAC9a97KLQ3XepnikchfCY4ROx6XljQW/w7Z13IrwbcKGln
QHv8ja5bzIICB3SCe3KCQo8FWoHW0ehIkYf9c6u11ygxXcNJeYP3NISkilIcSPx5NGLr9Dv6aNsKKpa1QaY2rCely39SNcPsFhMQHKOQsGZl6pnQWezGzSPNvUu/l13/
NxOy8/FeTh+XXRkPlltRH31FKE5fikB3n8aah826wa/xZgJA57cczZTtM6fnsWM89Rcc220qLBp4zlPu0RRUX/pVEfm5p8e6iDZ6DfM78LgDzUj32VlmfBOUxtFvJU5w
DmlC5SuGORuXNB46ezok/nVzWclE087CW6WrMnOpGN4efAw4Rl8k/1tWx7db2Y760gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mNSTRej+I45HK0oqC+8rtFu
xaqTkVM5haNmARDIXtLVMikNB0Qx3pFdWwwkj/6/SkRnckI1i/bOzDo7hjcWHXWnOZIOaATV5WaZ0+/AUfSa+hmnfw8FIwU8yBEqNgGa8eRKrgIUxO16DkclIN8ASv/o
/1o8T2wfswjjZ88jh3Vreb9tQ4yn3bzYzF3dZws4aOfDO90nz42ykyFM8HT2JYRDLqRk+Q/m4vIGnf19Y5W9O5GlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKU
OphwATLtaA5C0EoIoK1V9JkQrObRr5n9eXDGkf2vxdKHWZVFN1C4ZdsqpdxEhvEc/8OL8V/5n0T7YlGPctkvGsNOGTQdJtu7L9K4mRCRvGm02eVbDJxNS6yFi0AOzrLo
LXJ4OtesbURKs4dvr23SAXXAuhRiOcAASPBoIGAJnooBBVgWFnOlHtc8R5egWyFVdL/n6hSemlSoMGaUByUlc697KLQ3XepnikchfCY4ROx6XljQW/w7Z13IrwbcKGln
QHv8ja5bzIICB3SCe3KCQlmMBRKlyRoJTKQD7sGP/3SdqwDFx3Z7IeUKU7BdTFyyh1mVRTdQuGXbKqXcRIbxHP/Di/Ff+Z9E+2JRj3LZLxrDThk0HSbbuy/SuJkQkbxp
sgXNSCW7X6L/66iG8Syh+zRi6/Q7+mjbCiqWtUGmNqwnpct/UjXD7BYTEByjkLBmqKQ7xdDwFvvyXN54OdlDyyDLISLHgwIaGVLOoQjXGwoDzUj32VlmfBOUxtFvJU5w
DmlC5SuGORuXNB46ezok/nVzWclE087CW6WrMnOpGN6Wz0kh7fv3mfnJam44wlqZ0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mNSTRej+I45HK0oqC+8rtFu
Owk50N1RPlaKkvHOUr5dvykNB0Qx3pFdWwwkj/6/SkRnckI1i/bOzDo7hjcWHXWnOZIOaATV5WaZ0+/AUfSa+rC4cBpOYzDNXu71gJwtl7dKrgIUxO16DkclIN8ASv/o
/1o8T2wfswjjZ88jh3Vreb9tQ4yn3bzYzF3dZws4aOf50owVwigq8MWJgvkXHtUuh2ioRt3yDH9gq9WcbxqUqpGlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKU
OphwATLtaA5C0EoIoK1V9EMbTvYW1aSWG5GT7WZ4wzyHWZVFN1C4ZdsqpdxEhvEc/8OL8V/5n0T7YlGPctkvGsNOGTQdJtu7L9K4mRCRvGnmdxvgea207DubW/6u2Gv7
LXJ4OtesbURKs4dvr23SAXXAuhRiOcAASPBoIGAJnooBBVgWFnOlHtc8R5egWyFV3rrVtXY9dD1VmyWU57emioTFohwEY2DkMCTMZs86tZc9MI5bQvq0DRFT9Sp/3zYu
aY3SecHz2Z+yApnqIuEE+GbpryntX7HwLHo9PhKV0X5IPL8mMb6H1zueDkotuy9EStTi7MRKISN3e+5IDhyLV3XAuhRiOcAASPBoIGAJnooBBVgWFnOlHtc8R5egWyFV
gSiaIxEDuwVhqLCNY+x+5/6zTNgQ0rRvUD+LpVEG7fkk76a7Ht1Rj554TUjIMqWQqE9CrqyHZdKaroSYJ6A3VZb1g96bbH+1BTq2HuoIz6moJ7iTNMw/AAAzC6KpYw5Y
9zJH6MEfkXTWeH2tHzK6BT9jafvFoWcgzLH7EPp3R2KtG5/mT54mfrRn6WGa2XwxuHXNNsbrcONsfS09Lo+cvPnrmBBBc9BuX/FYWTvi6xpV0V0J9ZVXocsKnrBfI8ZH
cDaPRsBYw0KMX86Z0JTG0JqhPuIPr8wznqvpqTuklnhu1NyM5fwyusOGAHmWwwq8Fs3N1V02kZXkHoT+otXuhe+KAH3vD3WdC0E7QEb5ogLlbOPlYbypsz6UAmgAZjvS
bwiDpG2hf9xQjscjlqQ0Rm7z8jLJky8bT2ftqKhgcYkhPZuYVpydltCmziaeDv5DmxFTIkDtA5GNv2yW5jV69/7+mZjiBoliww8+DuRV3xjFAHj+iJOaeW9+xOLBrkR4
0TxzpJ0FCtCvme8DLmP/U5sRUyJA7QORjb9sluY1eve719hvOmk+eiQc2nFah8U2bvPyMsmTLxtPZ+2oqGBxiSvBj/hOA5h/lb4YSn1omWW6eIpeccOMFK5Kkim/FHXu
zxJ9zIYKZ3o4LsldtTOdQuSRjv0GsO4AXU3qKeON0Xln9kJ9PUoGZ+751Zl5GyM+Fww5MVSUZpPYs4sWiqlFdk9Y6CsuUC5kWDkR6JBIoCoXvAitdUkgp6b+fESH2t+Z
oMCjufuWjL57bkCI8xws7pYLLl8I/zdJGnvUYCkC09f4fjYkZhHCxEfgKXgc9KbhqNAOpARdApgYig2pdF7/3PFwiJ+SAGum/0tofiEs66VxU0NIHL16r5NXe09sJLq3
AzdEXZKcU57lFQO37kTQ93DNXNtsdT3bQzesxcDttgIG9Cm9GK/k7GDW+HHvsZn1xO+xRFZW92EgQqmK+3ROdApQmey/OPFV65E04c1foZVRa2LoyxFL5OeX6blHa4gc
sZ37Y8MGQpRUzXaaAxEe0u0tj2aeN8QUdJjBUqc3gqd+jqHL3Caz2KakTHYRUXa8soT2jBEeE8ypyx8QjmW5lVvp8Bj6VHV9OVF2AEMBWY+t5OhKD+R7pR/2VeJH54OD
qnHR2n4oKqVgGC4XIxNqprPHzb3DWVG5cVOnKm9RT3+Yd7nb05OOml55ZjGMO6XpCG+AGLTookLzCuAAN5I1BYb4D16clwRlTVs8/mlY7CmYvX8UWa+zzsDs9Mh11b8k
d/dbpVh75EdeTl41+3+aL3RnwU8Q1GwzzyePZy0cenKoSccfNTcJT7qLdpKsGOnDgKY3HOKtNh3t9dyzixdUhI47wU7vXAfKENEweIm0AeRWMHHxDst0YcDTSJm1YpPT
we0YZ6urZ6dBhSChuHZ0ZrRGtvWfjNgT0Mfl2Yc7LjrI5lam4UvfsoAoOMUpGUiUjjvBTu9cB8oQ0TB4ibQB5FYwcfEOy3RhwNNImbVik9N+uRNctBpDpWazL/O3u8f5
xQB4/oiTmnlvfsTiwa5EeDjNBCGPmDQ5T5zTzCFGaxI63Zu7ynaTpoQK3wQ6c0ipz79LXxpc7vddRYMkEsItnkQqacxCgMAZXIlmHd0fz/m+Lb9Mhd7X2ms6Wf3kytPy
uP2/D/RWtMivtdrkUos87rN3zIAv2NhTxYYTZSznLR7zLJup3x/2Z+xjdyymrXEEGjakeB0ZKPbrG+PJhpRJY8GmosDEPPccF/jzn2vca1wn9D6K1bYPpanW37xjmDS8
ywIrnOMTgk3yjeS2tj51p+PB04q5xjlfNNTd2D9Fs0wBOiaLivRq0H20uIOJWbehatFGxQF2nAZJHscVSOSCTRpFyYDcBRXZ29WxDYkdoiiZoD9mAnGxk+xk1TPK/Xf3
+B+NTxYIy2eDj3S3BU+ZqOl7Fj7STeyq34AF8+iUyUAwzTrMCwPa0nUafh2QBLA25I6HPuJ2ODEgKWjCRbifpBO+OlnH1kii5suV1ovfw2aDQhz8Vlt66PERuaha5WJP
RUO0n9T0QxkMcPrEDwZtvs6thaUv5jXHuWO0IV5xkWooPf12dVHsAbYkGRvZtbbzif1I1/kfvqZk2Ie394C41qgqI9LzgGnRVdtBsc6y6Ofsc2Fs84c5h1Cn+YbOn5RN
xTyg3jaOSa1rEqzarA/QfX1FKE5fikB3n8aah826wa/D7bkaZSjg31gI9RJjLKxUnwZtb9NSki9lvP6rAMZM8QPNSPfZWWZ8E5TG0W8lTnAOaULlK4Y5G5c0Hjp7OiT+
3E7/ssI3tWlbfPRO2YlSrIB8sxmUHlAqv9y4clzp7jP/quZ2O1gb9ksqyxwSuwFIW7z9J3VFbg6BYeC4mcQjyuUqcOzZ8Jwi/hp5e2SsZ5aveyi0N13qZ4pHIXwmOETs
el5Y0Fv8O2ddyK8G3ChpZx2CWqsMtBuqx//wKyhSXhncxVs4akxp+FvNxuHj9jEJ1kDeTQSet2EUifMY1sn83IukxsqkO6fI4SmyDiDPsGXaqSQH0rzJWmJSnR3JLNF8
1kDeTQSet2EUifMY1sn83AUH+dELbbSYQ0yHqM4MLyDIY+sK/WvsBLvwruMMYenzN8y/baK+7tZS52Ma6OfPzHXAuhRiOcAASPBoIGAJnorgszctdqDehH5sP/Wa+Pb9
XKqsgf48jV73zgykfxgT+DRi6/Q7+mjbCiqWtUGmNqz+4cAuvSY/V58BDExZGMNsFn6gkJaOa93APmvsvBjts6ulj06rOtMbdVH1RwKTctiet466qApO6GbyADyw6Fgh
8vU+RThaKAZgUNF8r72nd6ulj06rOtMbdVH1RwKTctiet466qApO6GbyADyw6FghrphHOrHbXy/Kk3SSJXDd9ZRIVVMAudvw7RBc+vEpIVG2nOzF9GBUAfQu9AJT9LHX
WM8YBGWA+D/f+MlxVQQbTimSi51MmhATA8bulqQ99xI9MI5bQvq0DRFT9Sp/3zYuJ78AR7LAQOx3rnlvExQ/bupt5fYFgXGhC/j93uCfMHGa4zOgIQhd48/t/+AOoH7w
fUUoTl+KQHefxpqHzbrBr+WCy1rjjIuVGCtMhJh/R4Dnh4lcLx1B7QEVaytGWcXZfUUoTl+KQHefxpqHzbrBr8PtuRplKODfWAj1EmMsrFSaMzIf89pa/PREZt9ZHTsj
juKysjij45Ilun990b45Gn1FKE5fikB3n8aah826wa/D7bkaZSjg31gI9RJjLKxUBVWqzecYaqgKQLPJqwVesZkvXbUmu2iJZwz6ytlJdMxnckI1i/bOzDo7hjcWHXWn
2YPBqGtfW5kk9tUQ9aDUVGFspv5IcoEZ08gzPSK1/m/aqSQH0rzJWmJSnR3JLNF81kDeTQSet2EUifMY1sn83AUH+dELbbSYQ0yHqM4MLyDnj5pQLKqgs6BhXQqQjjNx
3F2HRGMfwSi0qCI5lQmi6f3DkbC/vp3zYTAKcp47CuP7QCm3+jU2aael1QyaWw/kKK1inIdRsTckK3IGsYJMTzFdw0l5g/c0hKSKUhxI/Hk0Yuv0O/po2woqlrVBpjas
/uHALr0mP1efAQxMWRjDbBjTW0XQFxIPisnRbdN6EtVKrgIUxO16DkclIN8ASv/o/1o8T2wfswjjZ88jh3VreXkREfRRQE91LE3TJEGaEU2d25t7lTc7nAjjWduoZzfh
vGGmSNB4ezjwyuxCN1RxLYdZlUU3ULhl2yql3ESG8Ry6N+d/wtCY92VICekCyBqnmjHbxGkKN7mvzwN3QuDc79iirqSA6Bl4nMQ6WnHmkvr9w5Gwv76d82EwCnKeOwrj
+0Apt/o1NmmnpdUMmlsP5MM73SfPjbKTIUzwdPYlhEOLYSEnS5GIO0EJshHjU3iykaUI6BdDB4cBakAqvDTW0nHGz7FO4O7G3479t+2InFjDThk0HSbbuy/SuJkQkbxp
yNw8nno6iolko4R2xkebcH1FKE5fikB3n8aah826wa/D7bkaZSjg31gI9RJjLKxUCk1+Y6Vxga5grwEePdkXDx2eG+U5t3hW1UPPlIpTghfSBoqsTXZBfKS4CqWNm/17
wJ3dvzgrmwJcq6wjFyxiqjqYcAEy7WgOQtBKCKCtVfSaMzIf89pa/PREZt9ZHTsjjuKysjij45Ilun990b45Gn1FKE5fikB3n8aah826wa/D7bkaZSjg31gI9RJjLKxU
I7z16Gdp7gd8FyOwNOho4J2JZrIWCisdVRIxwCDaV1iHWZVFN1C4ZdsqpdxEhvEcujfnf8LQmPdlSAnpAsgap7qo4MVa0I9vRufFLah8e6wcM7FqWjavQFlSk9wQRShx
r3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWfnni2uiPG03BOTqTDCBQotceVqsO1D3xkp2l1edXJvG697KLQ3XepnikchfCY4ROx6XljQW/w7Z13IrwbcKGln
554trojxtNwTk6kwwgUKLek0oQcv2hu45G+umkUVjqkxXcNJeYP3NISkilIcSPx5NGLr9Dv6aNsKKpa1QaY2rP7hwC69Jj9XnwEMTFkYw2yjfsWuKq5lr+IihlDWJbcy
cdfjfrSy0VQIAlJopSs1nH1FKE5fikB3n8aah826wa/D7bkaZSjg31gI9RJjLKxUbBMkBLdarDzNcJvB4uvvHRSlRKD6e8kl2u2NNPrymXkDzUj32VlmfBOUxtFvJU5w
DmlC5SuGORuXNB46ezok/hq4cDkDBurTCac39dDl7NjBPL7pIzndmlXuAYyG+S/qr3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWfnni2uiPG03BOTqTDCBQot
zJWVgXUtNqZEKZVYeQ++6othISdLkYg7QQmyEeNTeLKRpQjoF0MHhwFqQCq8NNbSccbPsU7g7sbfjv237YicWMNOGTQdJtu7L9K4mRCRvGmOu0I8jwSItJcctk19aHH/
tpzsxfRgVAH0LvQCU/Sx11jPGARlgPg/3/jJcVUEG05maL5shwKiUv3ag3eIrkjLgbR74msJ17QOSRd+pmES4mJEjyFngoDu16siUxO8+RzEoSH0ygKLNmlOCfGIIYeI
Sq4CFMTteg5HJSDfAEr/6P9aPE9sH7MI42fPI4d1a3l5ERH0UUBPdSxN0yRBmhFNiEUPjDsssWg1Vt5Z7RbKONqpJAfSvMlaYlKdHcks0XzWQN5NBJ63YRSJ8xjWyfzc
BQf50QtttJhDTIeozgwvIK35tuZ2cDJhs/rmDp0NW3vdRtCmjxMu1Tk/rYLfeSkMPttlNocyNQ0I4jUrhX+1t5TZUjCPDpMWr1XXVnGRy7aYZzfYHTkVllCzG87DfQon
CEfuyt9rJtdUCHDmV0s6GjRi6/Q7+mjbCiqWtUGmNqz+4cAuvSY/V58BDExZGMNso37FriquZa/iIoZQ1iW3Mu5A6KQL6k8Sm0Dhs/y2WqCorqXdKFuVZY0h1osc8y5S
ZqRUs9KUdzslFr+p7PPCZtZA3k0EnrdhFInzGNbJ/NwFB/nRC220mENMh6jODC8grfm25nZwMmGz+uYOnQ1be3t575ZETWXfQgp2RWWzJ+AdcVRoF1w+oVewStREKQOM
MVoqVpalBCUENWKwJCQYg4dZlUU3ULhl2yql3ESG8Ry6N+d/wtCY92VICekCyBqnuqjgxVrQj29G58UtqHx7rEauZHjFsOYXv0U5W6CauX1hUqSvC6EjN+JM1BloexxE
waqghLKXV7SfxE4jDOvzRTnV5NyCT2qA7Q1ey2obC4cmdYcZQA5sVUP/q1wdi/zc7ZUujtwwhQ0cRlQa20J9KrS3bSl8aiq5Zb5I+aI33ItMTCBnDT2Cah/ovzKTc4zl
Ns+VYRj0vJjm8rcE4ogFB2pzh3pg94cKLK1vQ86njb3iU9a+AcTXdlExJSYiZN6GTmr8GcI1jgmpbVVTWDrqnWA0oOpkYO9thcHm5ap7/9xZfJb+rN79icRXi5mDupEB
SrzQMoVvSsmd2P+XdogErn0fn5OnZ7TAAp3S6LWtpVyxeB1aYBEhpzFZBeNRLDHJ/yAajXyGftAwWt+L+eIwFmDpvb7r68q35y41tG5ECgAEkjT0/SMaYb/MjE2fsdvC
VSHn0RFLrXTPvg8oVw9CKh86rjKkb8nghKApTXhTeQwctYQ6F8gkteTvZVGvJjUa+VXUyUcxSR8ojaVBMHs0Y6w4HGns5yTPlrVLa51nHdyDUAAQiCTO8BiCxIHnbG9j
GL8YNP3qOXXSIB4Rj+Nj7r+VCzpbfEAaFX7dYj9tmGY6TnrhdQHpMIOPU/Sy6mE7zREsQimt35Intlhs6t05C0lvTRegigbhy3a32fHRKvYlxWVmB0VVLnivOVJ4kSxJ
KnsLTsQGeDaOVZ81fGOxsN0qkfSLhsfy4Alj+lfN+MkXrfuddaD8OGMB4u1OrMgBK4yVlOyxA0OUPlA955Re51Om4Dtoc6VTO9IgwMUbG1s1QMi0b5mp98iSen2bnWWz
nH93K6kzqy+qj6qtgvi7xG0dJMul6zgeHMxKJ7hLkYrHUFPVUrZY2j800MxyjiV0bLHQf7AsEGvBCTmWSwjdA0SuqtFaC4ssy+ITOZpmGMdb/g2/A9DmxZjl22I4Pu4d
FRlCvkHB47nQd0yhR11j8W0dJMul6zgeHMxKJ7hLkYrHUFPVUrZY2j800MxyjiV0h5p0mjGEsgCHGyRLqK552FOm4Dtoc6VTO9IgwMUbG1s1QMi0b5mp98iSen2bnWWz
seZaIryvOTPbcU1TDp4FXH/hpoqEoKzZUrmj3ABtLTAAbbJrcyIIh/rwFzpZ6ELANLKoKlSL82Uu9oXjrBDzSFUC1pF3NxVDS5rxnsHYE7i/lQs6W3xAGhV+3WI/bZhm
zn2OuUsqQ+18bbCX2CVtJ0gZWxKtCiva2cj/JKdmxrZtHSTLpes4HhzMSie4S5GKTWMOn3Kl9EdNpVr1BOkwS1Om4Dtoc6VTO9IgwMUbG1vFKVePxJDExXR4y3mbCRQI
ZfNlJfMc1ur/IAYmW6OqNzWGj5U5eip5WBi7J9pnKulDDeD0j3FDeVGlN1qtpataOvXQaRm79iXCBXkt1cPsJqHxT4p+wISIoI8OT3P1GjdtHSTLpes4HhzMSie4S5GK
+w3TUwaLiA8nftIeaSCrys1oF948W0kqPUnLvgtw0dJTpuA7aHOlUzvSIMDFGxtbxSlXj8SQxMV0eMt5mwkUCLyAJlbaCENd2xijg8aRizoDaDsqqsfqVZ4tYtwPFVGh
Qw3g9I9xQ3lRpTdaraWrWuseC7xDflU0L3QfxnrfmGIVE50PFNojPvIbjqhsPFZ2SW9NF6CKBuHLdrfZ8dEq9lZ861sZbZEw/sr2kcOEVNOGdyNR3eJcdA6h7PTHYyS3
FtlldRlMJ6CEec1dQmMB+sWLmIJFAjV9f1zyAzuGJEa6IPPx6ALff05tmufLF9ooVQLWkXc3FUNLmvGewdgTuL+VCzpbfEAaFX7dYj9tmGa6e8pEiTCL+StpU1a5t2Wm
RzICF5AJTmPAhGnctoSU7ElvTRegigbhy3a32fHRKvZWfOtbGW2RMP7K9pHDhFTTHaFK4dbm8HpFbTsHc4pM7VOm4Dtoc6VTO9IgwMUbG1vFKVePxJDExXR4y3mbCRQI
6m3l9gWBcaEL+P3e4J8wced/USTzlZq6FvRSc7nk7vGOEfMyYXt5HPmQF3upyAS244TUZrp8lJRNZDKmLSNpzCTYb+tZ3g1PXzsRDGNawqltHSTLpes4HhzMSie4S5GK
+w3TUwaLiA8nftIeaSCrylwzLdqkxe4rddDWV954YSxTpuA7aHOlUzvSIMDFGxtbxSlXj8SQxMV0eMt5mwkUCGXzZSXzHNbq/yAGJlujqjejseuc3nJUjzsBaZRVKCIT
v5ULOlt8QBoVft1iP22YZlwfMgEA/ErLYpjcxwcpUWoVV9RbEXM+nZI+aZUsJ2kwQw3g9I9xQ3lRpTdaraWrWii0puaDV5vxMKCB1EoeC0faqSQH0rzJWmJSnR3JLNF8
htI/Vu8MJaYwqhb4WZAsFPYkYrONHeYqsSXreAo+AwNRPvD7lD6v1iO9pyse+DeDW/meqv/vHsqUxMV4jgKcUH/hpoqEoKzZUrmj3ABtLTDkqVWqT2053kVGjS/SxRXs
BVWqzecYaqgKQLPJqwVesfnHTtlOPHAbj6od2Y4fWjRtHSTLpes4HhzMSie4S5GK+w3TUwaLiA8nftIeaSCrym6C4X4mzphbxUizRg7nfigxXcNJeYP3NISkilIcSPx5
f+GmioSgrNlSuaPcAG0tMOSpVapPbTneRUaNL9LFFewFVarN5xhqqApAs8mrBV6xGL8YNP3qOXXSIB4Rj+Nj7r+VCzpbfEAaFX7dYj9tmGZF5+DX3VehRmaQMsOiRJSH
+6OweWkvwuWM6IY8GuraKCP8kAjBddi2uN9DZOUPGnHdKpH0i4bH8uAJY/pXzfjJA1AQuEYm69AATETrppRjcIqem0WwmGtjX1nRrSiLI1VErqrRWguLLMviEzmaZhjH
il611u1RgfZ3Zx42nEM8bDqYcAEy7WgOQtBKCKCtVfRBhBWNxW8Zp/BS6xWepWf/I/yQCMF12La430Nk5Q8acd0qkfSLhsfy4Alj+lfN+MkDUBC4Ribr0ABMROumlGNw
+ciZxQC5pMsZPbMG4ecguUSuqtFaC4ssy+ITOZpmGMeKXrXW7VGB9ndnHjacQzxsOphwATLtaA5C0EoIoK1V9NlrIU8l7qylQgg3+apMRxoj/JAIwXXYtrjfQ2TlDxpx
3SqR9IuGx/LgCWP6V834yQNQELhGJuvQAExE66aUY3CvMbd65iRBl/A+l59mNuUzRK6q0VoLiyzL4hM5mmYYx4petdbtUYH2d2ceNpxDPGw6mHABMu1oDkLQSgigrVX0
0+ORcIRuMLiA0STwwoYKtCP8kAjBddi2uN9DZOUPGnFTBmoWuZy0yJa+iGXEQZ9FjyqCMib3t6rUmTE+GHxQvMAKXX63Ck7+j7kx6Xx7Kx1pRp3qh8gVgwU4pknV+PsY
ZiZgHTPl2rJ2ojbsV7S+9d0bfdPZZOnfDpe596+zv6IEz7OH7NQB8S0bGD5jOdV74qJHZaPNRMG+vI8+0H8+UkqL6eb9UPyHPHho0lUh8eQTT3kBc+u1SaQWa4Woyc8K
8PUZrvwHxt2PNViA2nWv2ngDUmk473K/9VXcdeba0GlVAtaRdzcVQ0ua8Z7B2BO4nQjEVXnDrE1D1ELQ94lEwQhH7srfaybXVAhw5ldLOhp/4aaKhKCs2VK5o9wAbS0w
5KlVqk9tOd5FRo0v0sUV7Hqw5WD4a2vHiBeRYhxVnscxXcNJeYP3NISkilIcSPx51I7avMtgryDQY3vGHp32rB9hhH/y8PD+B/xl+PA+PCpJb00XoIoG4ct2t9nx0Sr2
VnzrWxltkTD+yvaRw4RU08NOGTQdJtu7L9K4mRCRvGnzoZ9gmIWvighZTQCUkL8wSnOYmHSXBqh+SIrEHsDpRtQUj+aCBLOtP2qoJQIY7yIyDZtaP39A0p3UxYI7LFAk
dW6Q1E9/cIXrO4pCRQAsAYnOfUtGzbrYemqP4y+46mSrm7Gk2lFFpKLWRcpfFmX9aEqvMnjwR2iVGsucp4+r75OumUaS+df6CwvjiaJDJN1kE3HOx9HGQ66FHRr2pWWW
6PIlKHdr7MTk25PtN9BYbQasYRFgXsgopH0fwgkWubnSBoqsTXZBfKS4CqWNm/17BobYEQ+Nh06EWNOfSwHiY4Nd69sQP5v0WZXttRuJ8ag3zL9tor7u1lLnYxro58/M
dcC6FGI5wABI8GggYAmeiiqwaiIQWSz4WqYYpV64rzSveyi0N13qZ4pHIXwmOETsel5Y0Fv8O2ddyK8G3ChpZ74mV+hKWabPZjO8ubL3Bf+19tSiZ0CJrMh9NPKW+Urn
16ZZIIeikEJe5zFDq/fSkbac7MX0YFQB9C70AlP0sddo/XMu18WpaxOLy37JDrN6fu55OAm8lsqdZbkMSX93kDFdw0l5g/c0hKSKUhxI/Hk0Yuv0O/po2woqlrVBpjas
J6XLf1I1w+wWExAco5CwZvpJvU9ytj0tFwCUDmM7LjoKa7Z0/ACZz4zA6ext4UYy/cORsL++nfNhMApynjsK41wyIZwcuUxMIfE7Xw7+GaZGSJt0EjPrwFS6PiVD84/Z
tpzsxfRgVAH0LvQCU/Sx12j9cy7XxalrE4vLfskOs3rUn10pSIsP0uCLFKRs0qPDDBph1c23vLR9lSbVAf3Bv/3DkbC/vp3zYTAKcp47CuMvs/pKtxdXMxWZHdbpncnE
54eJXC8dQe0BFWsrRlnF2X1FKE5fikB3n8aah826wa/xZgJA57cczZTtM6fnsWM8aMHT1JZT+iiqyE28wGZpvIJ1V1iXa5aaFj7eeJGC7RYOaULlK4Y5G5c0Hjp7OiT+
njG5+MjoHSBzabKA56oDR1yqrIH+PI1e984MpH8YE/g0Yuv0O/po2woqlrVBpjasJ6XLf1I1w+wWExAco5CwZnfOgR24GGMtunCvBhSCz/mrpY9OqzrTG3VR9UcCk3LY
nreOuqgKTuhm8gA8sOhYIf+2Wlkioek2vzHCj5gBWOmrpY9OqzrTG3VR9UcCk3LYnreOuqgKTuhm8gA8sOhYIdO6u3acVloCRG8UjuVrgbe2nJuvK1DvvCTiTCgt7hLR
PTCOW0L6tA0RU/Uqf982LmmN0nnB89mfsgKZ6iLhBPjVntmUynPQfdXuwDj5ovEz6ohZhz3Z2dxcYEtxdy668v3DkbC/vp3zYTAKcp47CuNcMiGcHLlMTCHxO18O/hmm
ml9JmquaRB4b5UE6n7UT2697KLQ3XepnikchfCY4ROx6XljQW/w7Z13IrwbcKGln9oII/VbALGvhLtE0xebiTv/rs720g1p6feJGrbWpXNX9w5Gwv76d82EwCnKeOwrj
XDIhnBy5TEwh8TtfDv4ZplYlXSq5GNHo+49darHUfz9QyAKw513dMclGvbcYkCtnel5Y0Fv8O2ddyK8G3ChpZ74mV+hKWabPZjO8ubL3Bf/rxXRzHEmuT21xASzshQKv
fUUoTl+KQHefxpqHzbrBr/FmAkDntxzNlO0zp+exYzztjxNWZl1pcRcRJ50RIZKWq6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCEpuJlwt9rvEBNqDQlLMAdo
r3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWdRj2cPeJtfxjzHjncXQNBHH3pYHeGIMVjuvBnXydBB79IGiqxNdkF8pLgKpY2b/XsGhtgRD42HToRY059LAeJj
oOalr/oGi0N8MzrqLTGbMOfEJImKdfu0J54BKa2crkB1wLoUYjnAAEjwaCBgCZ6KAQVYFhZzpR7XPEeXoFshVU1wrDqGDbGOPzNsWeahryjSBoqsTXZBfKS4CqWNm/17
BobYEQ+Nh06EWNOfSwHiY/bbpLSUqU57dPlnQ9ysqJ2rpY9OqzrTG3VR9UcCk3LYnreOuqgKTuhm8gA8sOhYIdO6u3acVloCRG8UjuVrgbeOcmtq2PzIpKZ/uP+O9ljL
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mOg5qWv+gaLQ3wzOuotMZsw58QkiYp1+7QnngEprZyuQHXAuhRiOcAASPBoIGAJnooBBVgWFnOlHtc8R5egWyFV
sJvRGQM5E1elN5u6Aw7bhj0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4QEuYZk/UBt/RUFh2GoPRbAPNSPfZWWZ8E5TG0W8lTnAOaULlK4Y5G5c0Hjp7OiT+
M6Z2gB/d5bO4DGWjQyfri+rYw+n1SBpI0PcTstXTXaU9MI5bQvq0DRFT9Sp/3zYuaY3SecHz2Z+yApnqIuEE+NWe2ZTKc9B91e7AOPmi8TPqiFmHPdnZ3FxgS3F3Lrry
/cORsL++nfNhMApynjsK41wyIZwcuUxMIfE7Xw7+Gaards7rQN4KOg/DEiekbe40PTCOW0L6tA0RU/Uqf982LmmN0nnB89mfsgKZ6iLhBPiUbZkDCkZ60EdxWTf4d7E2
r3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWdRj2cPeJtfxjzHjncXQNBH2qm0R6dvRZLhS0o+i80YCz0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4
1Z7ZlMpz0H3V7sA4+aLxM+qIWYc92dncXGBLcXcuuvL9w5Gwv76d82EwCnKeOwrjXDIhnBy5TEwh8TtfDv4Zpk6j7sD0gEjBF6XWhbblM2erpY9OqzrTG3VR9UcCk3LY
nreOuqgKTuhm8gA8sOhYIQEDUZLKoHq9X5VBfEcU3LixlwwrQM82ZnZkV97EIDgX/1o8T2wfswjjZ88jh3Vreb9tQ4yn3bzYzF3dZws4aOfUIAXi5t1FtyoJgotx79cx
PTCOW0L6tA0RU/Uqf982LmmN0nnB89mfsgKZ6iLhBPjVntmUynPQfdXuwDj5ovEz6ohZhz3Z2dxcYEtxdy668v3DkbC/vp3zYTAKcp47CuNcMiGcHLlMTCHxO18O/hmm
z5spKBxr7bQAO8PLLZB4xNIGiqxNdkF8pLgKpY2b/XsGhtgRD42HToRY059LAeJjgqOSnxVbbWwPWdcC0ThojD0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4
JyIU0B8hrSosy+pP6V50WwBdgb0Poa+TPpRNYNh2k2KRpQjoF0MHhwFqQCq8NNbSys5+d1LWLIUzk8A4UjJClEtllc+Gk1ROzrnyQP1EXEaxf/lovI4iZIEXxqqYxC5G
DmlC5SuGORuXNB46ezok/p4xufjI6B0gc2mygOeqA0cOzNZacwQm+Iu1NCnFHOSPkaUI6BdDB4cBakAqvDTW0srOfndS1iyFM5PAOFIyQpR0haQ1nLg6FKqgxKahkj02
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mOumEc6sdtfL8qTdJIlcN31+Ft0HOtD01sP3a6RJXJ2YJGlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKU
S2WVz4aTVE7OufJA/URcRrF/+Wi8jiJkgRfGqpjELkYOaULlK4Y5G5c0Hjp7OiT+njG5+MjoHSBzabKA56oDR7krOMN72XLF9GZprmyhsw3/quZ2O1gb9ksqyxwSuwFI
SNZodRTQofIbQ4VJyf6YGYEkO03zka7dB4mgBIYoIi1D7DTU4kl8qHU3ktAHrrzYsxBfQTbqDNodXE8XP522XencajSB5R9DBo3qqRtAYym4qrQZDcwWujDcuwR+FUoV
n7RIhfJtaQTs7dnMnWqdlMD+IiR8XaCKl6MQiA19t9Ph8K9Y18y/7MjfDkscE6gmHTdAJWZY5WJrWQ6+qQ7UyzgMrH9Vw2Tc2zp2zxRRBATzLJup3x/2Z+xjdyymrXEE
7vhjQ8XTcSg3fwusAA6zmWfQQS9nOKO9YUJEtuS++XYYpteFhLq+mWRculJKOowJnYYIs6sHQWSy63i+1Xf6v/6rA3cHMP3pDAibLLfsgGSm+gqBn3T6R7CpvC/fo/kp
E746WcfWSKLmy5XWi9/DZm2zClvWldWxbE/ZFhDrWrMKyFYTJpP0RnUcwrnUnDvd8dOkQ/xXyLq+W/W4oVYgfmFSTUDntpfbAjJanlpEXb/u+GNDxdNxKDd/C6wADrOZ
Z9BBL2c4o71hQkS25L75dhn/wxWElJHHjYq7i9XTW8dT6LMqle0aIPkXVcpA2ZJPhmC6QV7FBNuqpmzxt7OOYVvl4kQ/f9grxWTHvaDqyWNm/64/Ch1sitprKBWwMqzB
k/vvC/jYRT12so03ToIbF7oyquy2+YsYeXBvirbGNgvyilfU5Jnu5AhTLarAciuMuP2/D/RWtMivtdrkUos87moFHXu1ZCmG3bhV3wbEcCHCtnWMrcRIBZT64bi1Ap3r
ufqm4n/adSWBiATP9D3XIRMIY05zkh/ThAOMa3wD+ZW4/b8P9Fa0yK+12uRSizzuYbFsC1xwKDW8mIpaSoWTZZP77wv42EU9drKNN06CGxdhFvMjZAIYRjUP6qbaWioJ
5fG4ZRe4e5fOmuAthb8huW3DnaH99wGILBQvHfpyEY9lL14oNYYl8oQ4/eLCFWb4VO+f4kOVE4i3unKTwt+z9oOpiBDjkNCGEwJJDjihocZNjmGYdpLz8gY28yP33LOH
gOs3ZMoNVi7rykFFzK8heL+N842JrSosXhY4rw4R7UacEvy2/rP5JSYpkJL76KL0lseY0QwoUqNoPx1OpoNSrB6toZGU9XrdQSNJoHUUQJPTkLpeemU3UBWNX1HqtqZO
jsNmP+FUPex9UHdcEAnf8cOeqKMJ2S5uKAbKhfAm1FYJ7P22RFhhrIxhxKFTh2yC7d2TH+7JQB644b69n3wSGR97aqGs86folIxfsdZemaiK8gYWmQJb/r0JFD7reSQl
rZAVMJhttom2tDl6Mt0nTTa5zmDY57Uf/npYSekQ2dmyQLjaUdt2/zonnz3m3FbMXsRYS+QJL5ncUPlXBY3+f32WHAJpYtsb19lw1oo+aGgAx3GkfaF4NFGkpwHBBsNh
jEsF9BOsBJdta54FyZvg8O/mu9d3l340UuqZ7x0lsZFE/YzMIhY71ze0Fs3YRxmpYtkSFpHWmUPN9F8o8AN7KsI6zTeE35BDq0oeKIydoMvO+WSuEazdF2wIzgboayUU
r2Oja9OH5WteH1G+nrZlqXnxSRMJm09Dd6A+rBsv0EqFCLD6nA6Hp5gvlGIkA4AMnt7DcE8fmgwP06XOkaoSfxqaXf25NW/q1ffSVL+0C7/972o+/kdgA36cYmyOyGu1
SiI5jtxYyncWj2ZxguMZz7vcLrfHSCF+iPZdUMaRGrRRr+qNDmK5bkzfvsFeMNYnrZAVMJhttom2tDl6Mt0nTTk5eTLEg2GNphNUI+ilb29nW5aElwXZK1ZgqUdOJPkW
u9wut8dIIX6I9l1QxpEatIYkETdw+g3bdwEuFesRcI2tkBUwmG22iba0OXoy3SdNxQfY3zHaKAkt3wNwQ6O0vppsx2NPk2R0X62K6EUiWpe73C63x0ghfoj2XVDGkRq0
KvuS4GRlghnSMGJu1+zPWRsgGucsw3WPoDYg3UN4RHzT/QlWbTbsaIHkcd/f7edx9pM1ylRquX+TqSurMrgogduZrzfaYCC6o2I4WuFYc+BLSLmXnhzWTUESQLkTP6uc
B/u8xndCMEuXOiuwLT16R+R0qEeww6ir/UFeBh+C2+QldQe4RVVDIeudhlA/YbhSXDeubRbkdV/MhVpmbQjSpj+8CluYsFXcUtamgYIcmDLvbwkpS+n+/TGH+IMIrNHL
NjbbUXnnV3WcsX+Ui5h74GRcY4m5SnaXKi8N1BMD8VThW4+vxZh5VxqDl8ApyGpFpETu9tvDDkZZlT14AvqHMqBHw0oHVbnSOnMuhJnypSKTlGk/ikbd1m/8KmQPmEAt
GxBhar7BJwOJTut71zEW4+y3GsV8Wn3kxq7WezeErO6wgDCu8QvMj/tOzQ5Y/eMgOAJ7fu5k5nZiSU1aUuR78/2uDHkpOale2io7Ypr9Of+G+A9enJcEZU1bPP5pWOwp
2NqKDxsfnUQt1JNmzThtzKyXnT4K4tp54r64T8ICybYjK8mVNlN7y0QAFuOVw2Bh/7aclqenp62No5Ykl16XoXvn2wF2sWfYlh6bGHG7pp6JkMcw2GkBC8u2ivsVsv/O
LIFy8o53AwiXW0ielKcE/BNABH2JybuqMVJZnQUQ+MQ+vaLl7ZGc2mJ2PAMnmKl5mazWv2lAWF686LMKXwRf2aVGcNwnhgLwJit71XmZ+7dqR2w+Kd5iEqpwZ3N6fcmu
soeGE5oOhOgxydHOyCwNtwdjSk1plWACFrpAd+XYp1hxAWxSccJa8uxt/PkM3rbEK0dc0jyfeI2C7kjoE650jroyquy2+YsYeXBvirbGNgtNdoioUAHy0IH53yL48MHE
hvgPXpyXBGVNWzz+aVjsKVHozByeernJPVQCB6rFNRX7HBl5rGQ9MZJnOLDBRZuqy4ucOVJdP1qgObTAZcYBa/1DG7pwHRyqCPzjd/6r/VTWQN5NBJ63YRSJ8xjWyfzc
n6idFNTjcyGdFocxjFlNsmZovmyHAqJS/dqDd4iuSMtwqMaO1oL0f4uU6rPZhieATQgpui1kSkD09TMlH3otgxSWVdnJg3GoMEueWFIEHRiRpQjoF0MHhwFqQCq8NNbS
ys5+d1LWLIUzk8A4UjJClDqYcAEy7WgOQtBKCKCtVfQpOcjoAh+OYrDvcPzrozzUW9QMhXWvXDtU+RWN5H29YsDUuStATuFGdUJx5/R9cpuveyi0N13qZ4pHIXwmOETs
el5Y0Fv8O2ddyK8G3ChpZ0B7/I2uW8yCAgd0gntygkJX2eP13UX/OChHCWeI846KhdzP0taeNftozUVdf3+VwafX8jghJY2KiMFhN+T/UkzbAxJSyla9AsypGfJoa7rw
fUUoTl+KQHefxpqHzbrBr/FmAkDntxzNlO0zp+exYzyt+bbmdnAyYbP65g6dDVt7PhiXU5biy6Xwi3mlVcQ8Q6iupd0oW5VljSHWixzzLlKz0vY7+n+XG7+lohsA7eso
tpzsxfRgVAH0LvQCU/Sx12j9cy7XxalrE4vLfskOs3pAt9w3BZXKqVM8UkrHqlw5ySFRV2FohWo7iM2unSKjX5QSCB0YesozkY+PO+tqKdXfMLtXBlRPALLv3qit1rnJ
r3sotDdd6meKRyF8JjhE7HpeWNBb/DtnXcivBtwoaWdAe/yNrlvMggIHdIJ7coJCORTAgUUiEEgJlMyNzqjfvdqpJAfSvMlaYlKdHcks0XwwLYIvgUlACVkSTGl+aFUx
TCE288DkFHI2wsNNJN2m2n1FKE5fikB3n8aah826wa/xZgJA57cczZTtM6fnsWM8rfm25nZwMmGz+uYOnQ1be7PR3uURSNWzbzcV8PIfbtodcVRoF1w+oVewStREKQOM
DgBSp5xHVpmaK4mDWun1Vv+q5nY7WBv2SyrLHBK7AUhI1mh1FNCh8htDhUnJ/pgZsuGgY4ulq2aX2YKDLM1hI9O4newRnp9wDmfmYufrDalgB5KcQCC/dxXxZCdAFEht
AYQtVHyaZ5bzrLk3nib4gh34X3Xk8fWjaj7a112P+vwOaULlK4Y5G5c0Hjp7OiT+dXNZyUTTzsJbpasyc6kY3rBB5//ZPlnlbALBI9WK4wUxXcNJeYP3NISkilIcSPx5
UaW4fX2pBEJnZuYqxpkCabEz6EBbAuMpYmaU+kRXlApnckI1i/bOzDo7hjcWHXWnOZIOaATV5WaZ0+/AUfSa+qN+xa4qrmWv4iKGUNYltzJOxmOAS2+qmzlptFUX4UBW
qK6l3ShblWWNIdaLHPMuUtKUhDTHN33Vn6Scdj1FkyeRpQjoF0MHhwFqQCq8NNbSys5+d1LWLIUzk8A4UjJClDqYcAEy7WgOQtBKCKCtVfR4dKrYQaaTo1tUADnJNCZA
LXJ4OtesbURKs4dvr23SAXXAuhRiOcAASPBoIGAJnopjgE7mScx4A+w3mCj0Wm/tSizFUMMSLgHE72ajbHxFLTRi6/Q7+mjbCiqWtUGmNqwi2EpQUtX+XzFUyQfBsDb/
h+BsHMDklstj3l8YBReCWP9aPE9sH7MI42fPI4d1a3nTmrTDEy8EFSlKb2ryr7I2RCasRiekg0qNSy0Jy+/uckNWjtWM0p4DCxUBQGjzAr3vsXcp4Px//J5yqdDtLBXF
T9qhYUh4EG8cR6duqR+f9aDBg3DxOIl0JQw4HA1nEZ42lK04+8oNmLzKCH5ebIif2RlnH/LBliaNK8XLrRCMl75nFTHcLXEiOo+yxf1vfZgakAT8yMIf3e6OlE3qU49W
UO09Rf55jNDMqKBuPkule8nYgNKLLnCPob7uZETXRNgL92stq1wIumRCqzbC5NWIPdy66MGwjpliRTpNvHjYJd+aykyWYdbxfskZvDrPSs3Pm1dTsJ4khPpRJfLGaGZa
7IxTf6T5elHYFbJj+vhhuQ6AoIFPqeiH4LJ2z3X2xP9vvm3rwLddSTaMxeSPDafoJPh677B2YLRwYWFiUQpraJrNY96LxDxbKknZohg0rE9B4iGLqOGeADLjbOhjieS4
Vjo/kA2REOsbp41a2hVhe00IKbotZEpA9PUzJR96LYMAJCIZJ24Ql+g80CsTBoGts4+auKDpDRaaAlDwlnNoYrUsGBE6uieesor/W+WTUipgB5KcQCC/dxXxZCdAFEht
+AcXZzxOoCAfFIN1eBeF4lkJuipZ3qqtHYkHQmSKD3vDLKIn41HXy5tepFYIHHS4f1RkxobQWgg1pirkN+g38NqpJAfSvMlaYlKdHcks0XzZBphb3tbncJ6rN9QCoSuD
WONW7gH0crsnLdiA328VcbOPmrig6Q0WmgJQ8JZzaGIhJZx2hSlwc6oH0byyieFj+RPug31UuHibMStN4gjZZ/MskxaJufkU2PtMup8JrNeDucgmMSdCKZxg6ZEXrl1f
zUBH0P+b2ClmLFB+Gv9Cs7SplEXPojD85fFpGOu8xBtb1AyFda9cO1T5FY3kfb1ieC6l8870erjZ3rMlgD5kUbOPmrig6Q0WmgJQ8JZzaGLnW4nehkeajE08bzRzTeVz
peufOAyMFHTOvyxtg4QMzsKhSfxzULkeH5XTuMaa95rPKMcMYavSG+ZiiBu9iD/bkEjYo2HFJBNlbQ/xQyxIPTR6JaRXRc47QiNYw+CIZ1ioB0sUjm3tHzUn39Hk67Fd
sxDjj306QZZNtMgPs/SuSilD3JtqOpFVrL2SRlaIvqnfqvrvXqgR0nE9VotiNodQIi5k0S84V6ZS8qOAXMN5Vd6uoOZK+Z9A5qPJ07kQKjo+2tfwBUhzE7eHUxAahj//
XgGAu/PnkKgNWe3IqOmHSBxy8Cs5NQt0XdEKwZE5vUdzwNMR111dv4gyZei8uS1O42qgGdGrjQCBTslgJxRF+E0IKbotZEpA9PUzJR96LYM3TRgeVYBHJ22T4IYEOvzI
TQgpui1kSkD09TMlH3otg4Loh71x4qsHFWAB5wpOXsggMNPxcdu2T2ZxOuHcZH4WHXFUaBdcPqFXsErURCkDjBDmepKsyEgsijzhlaAlN/Lbcf/niNVgoz/uxoNTy/o2
HCbwIb9tMK73zoatBAt0heUqcOzZ8Jwi/hp5e2SsZ5Zb1AyFda9cO1T5FY3kfb1ij3d9D3UXozMAstxgm1GiJ/E822Nv3mCN8IiK9kI9FsjDo0JfxhN5McUnMcwEVShU
VsYdKdsYb8ZnnCqC8g+xg0/4E0MfuUZRLR9sf35QWkwnjJroaNF8zOJHdm1dVDaJO76S0FP1Y9mORCGN30t4FzNMfAJ9ZEbjTyYJY/QJXlOPd30PdRejMwCy3GCbUaIn
XKqsgf48jV73zgykfxgT+MXGi3hrgSHOj//GBoZjspwjj/BKhTa47wYhUkLt6bsdn5CzHCPB3JbjnjfV1LBZ2iNLzCHyCltKYTUwz7TL2ig8bKjn3WAEld0r7gb2OicL
HXFUaBdcPqFXsErURCkDjGu9wl22W+9Bi/Co64QZgpFhhH2mZ3xrTDtiCpdYJ0d9W9QMhXWvXDtU+RWN5H29YoaImTht+0P5xFj1ZBh5OAGF3aRqhzqDZZ7BhlBgKe5s
66PGK3Fsg5oOtpi8O8a6mSeMmuho0XzM4kd2bV1UNolhbKb+SHKBGdPIMz0itf5v2qkkB9K8yVpiUp0dySzRfN4jqlBgIBV7GS2Pry54y03DThk0HSbbuy/SuJkQkbxp
LsdeJ/yaAvikmxB9uXW2HsXGi3hrgSHOj//GBoZjspxKi+nm/VD8hzx4aNJVIfHkW5t70yyFQycNHPzxpcNX+B1xVGgXXD6hV7BK1EQpA4wRA15PQANfOAEf5hJKUSA6
qNj6iPEiMCh8wCI14HaSIBwm8CG/bTCu986GrQQLdIVAt9w3BZXKqVM8UkrHqlw5zCwaj9lUYH0u6hLOBU5hJJQSCB0YesozkY+PO+tqKdUbFt9dq8c6ReF+d+oc7ZMq
Qg87++JbycVDtajDF2CkGE0IKbotZEpA9PUzJR96LYN72XigU3os0LOR/8JhPjqQ1QotJShNGedyyvsWEWXwQT4C0VsbxtJqOftlQc0rCHUcJvAhv20wrvfOhq0EC3SF
QLfcNwWVyqlTPFJKx6pcOd1G0KaPEy7VOT+tgt95KQzWQN5NBJ63YRSJ8xjWyfzc1aN4TXcq8iYXu7plxrx41dqpJAfSvMlaYlKdHcks0XwlI6qYd+rj/TWvy4kIMMBH
iF3UV5DTuZoR+CizNeJtvk0IKbotZEpA9PUzJR96LYOfwVP6Mi3hp/dAduiYU4bDHXFUaBdcPqFXsErURCkDjCu55RCbptIu7WVPHXuy6t9GxlLTeKBcuFPdV/mysyN6
8yyTFom5+RTY+0y6nwms1zgfgzY7QfdrEFvpBmXASoPzLJMWibn5FNj7TLqfCazXZfNlJfMc1ur/IAYmW6OqN+B3Qk7fxIOZyX8lOy/e1u1X/Yr4Ly7ww+MbVhLn8Pt5
d953cPLFOudctgb30apQmlf9ivgvLvDD4xtWEufw+3mASm08k5SDYyqSDkd/mQb4PHdFGYdX5RIiT2sVV5xHCRsUJ7cL8altpO7xMoEUD50+PeYNdn1GZDYubdJzzlVG
eeaofWixv60vDrnh9shfQ5AkM4sVgj6IjptTWnELMggFTNf+juK880vz8jdPp0NwvA/h+qbkAW6jq7KBXh2VZ9EmrlcfzPnmrS3uLr3EYR9YXyTDiQ0Cb1Ftw7c/sLpn
3VTeT6s717Xl7j1Uwpwj4MG3WHQY7gX/+bgAlWHDAKTyjJW1LO7jz58iHa8T+2cJeeaofWixv60vDrnh9shfQx2T2VfwfCwLD3J0SwEzHSBQU7JPwDMX9OmXT/WwpdVc
XxhULNHYXaoR/kCmXPnSUgVM1/6O4rzzS/PyN0+nQ3AraEX5hWn3HLHINJ/vzssV2Vir1qCck0ZEEkXieQ1SzVxSXg0jjJFHnwAHXIi05Un9v2y+fmY8m6BgKu8QuKBF
v+TnZzKxiZGKq6R0TUkR/+y5rsmsOnVyW00N86vHUXRQU7JPwDMX9OmXT/WwpdVc+HhpKoKPWnlKBcwYcaNS/psgONPYbhoTSBsJYYf0xjPhHPFFv6Ijc+fmJdbJPWWG
jfAJ+AjWzeT3Qxpi3IduVtEmrlcfzPnmrS3uLr3EYR/i7e5bvtLrG5zFiVbm6AVuV/2K+C8u8MPjG1YS5/D7eRStF0Dmso/emAINisMFZVSTNlCZubr32O7ec52B4xvW
zgXJLl1floqTir//hwXhTD0iE3aBf2Wtg4vaRpERURJ55qh9aLG/rS8OueH2yF9DxgFv/55Fh674ao3Uo/CTQDF7fDtfaNwlKMLTD5ihicLTb0XeWXEjGnBH+MHmM4Tm
f2eA1mRJJJZY755xRuamETAWXvCZhPB7GCSX+07SOpgeGbE0/vcLjlfaMFE+QZKxv+TnZzKxiZGKq6R0TUkR/9dfMOV8hyi+JQTozerVI0eDMJXs+7m8IRpdzfVUHKFd
hPN1b9aH9pSYs+uasXSbfEJUvtt8NEacnrL90ZW0dwdFx9X836xgjd0lrWlm3BGYeeaofWixv60vDrnh9shfQ0FvnXGrpSa2G0IL0mXvA3SUEggdGHrKM5GPjzvrainV
9s8oW7v03dmaaynex41gDnEsmSKomv7x+st1ludsXeRNCCm6LWRKQPT1MyUfei2DDRy3pGCn+TwyKehKzuXTUmft+S7InqX4oGYklAastQWu7BYmW3z4YGc+FokUft67
8yZpPXKFt2LmscbUnmKGCPwNIn9Kc0YHIpXlUc1IBOWDkSGuYaqOYoNIjN7WlFZuYAeSnEAgv3cV8WQnQBRIbUHdgbK+zP160x6kSbSiy3WrYgCACxxj3DOVEitNoEit
M0x8An1kRuNPJglj9AleU5YDJ3UzgayP4irPgnqKR4pcqqyB/jyNXvfODKR/GBP4/vGWjfFLXZkkXEggzHcsbRHEL6iR9TaCMn6EUcVacT9b1AyFda9cO1T5FY3kfb1i
Y5zDG8c7nNDDozCUh5V6i5QSCB0YesozkY+PO+tqKdX2zyhbu/Td2ZprKd7HjWAONWNJFLQ45g4IKGaK353sWk0IKbotZEpA9PUzJR96LYMNHLekYKf5PDIp6ErO5dNS
Z+35LsiepfigZiSUBqy1Ba7sFiZbfPhgZz4WiRR+3rsdnoa122opxcbVs/vgfkH8/A0if0pzRgcileVRzUgE5cM/nPOsHhgoWR54w7U6n1RgB5KcQCC/dxXxZCdAFEht
Qd2Bsr7M/XrTHqRJtKLLdQC8kDxo5nUfLwBUhRJeDMR21Eo16bnR/tx7jDV/IhM0GbEKAdFtuztr2Ylf51jKzZbQU4T5yeYB4VRMWLgs3C72DAeHqCM8yUaoIdTwJRMR
ZXwoFrakmWkX6MLIa5BzUd+2cNMk8rmQSlStC53i5HOYQxcdFdQDjUxuD2EcQ4fgMV3DSXmD9zSEpIpSHEj8ef7xlo3xS12ZJFxIIMx3LG1ATSCZ9i73mT+nKtizQSUL
cqzVscU9kfWX/NCSXL+XFiIuZNEvOFemUvKjgFzDeVU6mHABMu1oDkLQSgigrVX00sKEUTbuMV8fEdIY5ZP6V6iupd0oW5VljSHWixzzLlK32jVw8+q6jSyf0GXvz2a5
2iNxFDmxzeHhbPj7+zPipk/4E0MfuUZRLR9sf35QWkwZsQoB0W27O2vZiV/nWMrNla2u0WJCVd726sCoHVnbAgg5R28Z3CCX4uQclfmVx//2zyhbu/Td2ZprKd7HjWAO
KK1inIdRsTckK3IGsYJMTzFdw0l5g/c0hKSKUhxI/Hn+8ZaN8UtdmSRcSCDMdyxtZmi+bIcColL92oN3iK5Iy87QKDCoDcBcjNOsbC9Q9VzXKiLN0Kh45X8Ab80UiH/q
9Rcc220qLBp4zlPu0RRUXzbOs5QrL6rQhFstBxLCwftNCCm6LWRKQPT1MyUfei2DeJ1LUFLI5oWSK53dzEDlwG7NeNzerGGad8k6QRBhIl/zLJMWibn5FNj7TLqfCazX
suGgY4ulq2aX2YKDLM1hIzezwmiyOHEY4SC974MLXnKl6584DIwUdM6/LG2DhAzO84izBkWoasb4tovD++gOSayMWKevc5JLdCrZpeKh5rsIOUdvGdwgl+LkHJX5lcf/
9s8oW7v03dmaaynex41gDjPxvQbCq8IUxdCPupYqSUP5E+6DfVS4eJsxK03iCNln8yyTFom5+RTY+0y6nwms17LhoGOLpatml9mCgyzNYSM9vC2bDk82XnDFlVar1IGP
9gwHh6gjPMlGqCHU8CUTEUC33DcFlcqpUzxSSseqXDlCqIF9JCNtGjZ+/myzgbY0peufOAyMFHTOvyxtg4QMzvOIswZFqGrG+LaLw/voDkns+ojsJeceojG+CHP3v6jK
Sq4CFMTteg5HJSDfAEr/6P9aPE9sH7MI42fPI4d1a3mmaMvF4VMtJdYplmwaAySPT/gTQx+5RlEtH2x/flBaTLCjRM3nJJRAVrzWnArGeHSdmBRDlCJS+uTCFnogWs6a
0B1H6V7DM18gb/5kgMBdpxNPdyIR/8FtJEfN8jPmpYXRJq5XH8z55q0t7i69xGEf5POTGetjR9RqcmU/UZenDUlvTRegigbhy3a32fHRKvb1HQsNl3vOn6rWAYxIi+Ui
62nY+jShQU1XLoE9PSsnYlhn7rca2mmehrW9BM2crGxLaMmw4q7rjC+dorsgGiCbWGfutxraaZ6Gtb0EzZysbIRyvXa+Kzq2PDkUx3yY1bTZWKvWoJyTRkQSReJ5DVLN
LQLOHcaHA0CRE7tT+iAeECA48VxdviCrBUfSwxvqejarnSp0hxRZ6IDmPrCmWnxaLKngFR7CA6IL3LKKesW5b9Ev6g7+wvIm5G0OXmBBYga3b/wvYJ5i5vMaVFPIEWn1
MMf1VEOdABUddtfV9UGxln3UOtTksuq/SxU/hPBLz308d0UZh1flEiJPaxVXnEcJltH1GOWSY8vyZ2v6qDEC6urG9vmun3/OdxqH2e8eWWernSp0hxRZ6IDmPrCmWnxa
8Sd7TwUF8NWIKiHhOBE09dev/W6FdlrGdKlWKtO3eeQGxFxEKL369BZ365/fGgBB48ZZNj7V0jfQ1HbfrXjHFa6Sh3g3kU2qO96BLbLeKwWJlV+8IPBEVlwE4bA8pDFU
T1grOIBtZbVruCapn1gr124w0ICRxeorulT6UKYMA8Y2UOtyVY2zRYHSzPRD/6pNTz1cNO8FtZ2lfI5iTsZo0dev/W6FdlrGdKlWKtO3eeSUjHqki5pNChElyswYRDBR
9LbtzDyN/FS5BcqCEYDPojl/FmQitsOgkCdMyUoCiSOlEIfXONwF4nwOVf98LodNMMf1VEOdABUddtfV9UGxlt+xI+G0hm05bdTYTpnr8nVYZ+63Gtppnoa1vQTNnKxs
beYGJUCi66ZTy/2IxMEUVR4ZsTT+9wuOV9owUT5BkrGrnSp0hxRZ6IDmPrCmWnxaiHJ1xZrygiVUNwZ0mT91x6udKnSHFFnogOY+sKZafFrnsA/1EruMLu+AFOX+6wO2
pG6BclAttpcVcUBfbWlEswIEVftCt8J1u0K9G2CnK2PPUEhHr6oyAMRiM/p5bl7kybw8Kn1T+I0RUq1bYIWL7s4SEdKPaPsN0XmBfbeZamY2UOtyVY2zRYHSzPRD/6pN
uqEXJvB+3Fo/I/JV2rjjbC0Czh3GhwNAkRO7U/ogHhBUHTDf7MhViZJn+Kue4P+efKPFN7oPYkwcB1rtTCsNJBPSkaQT4P8N9dlXUKj7kMGrnSp0hxRZ6IDmPrCmWnxa
gPnGh13xdUrNSehvTR9Ph/mE0/THssovMK3o/4oSz9nFi5iCRQI1fX9c8gM7hiRGANaT3UrjH+eKms2CprWhGOPTx8hFBvRrvQrHgS9TqueJRCUYAHThVdu53iUlDy+0
5yIM9OdllrMKvacu7WJvC+FzcmBY5eLreHNcckBJcsCNzkfsDmGKZilVgnioovMymhkanFoPXUDPSK+P1pYkciTYb+tZ3g1PXzsRDGNawqltHSTLpes4HhzMSie4S5GK
slQbHSJn7gGH/HLjFd4NWAoUJV2L327STRqBuyXZnZXFXeSGmDWkt2iWwF/WSGNjQw3g9I9xQ3lRpTdaraWrWthtMR/4mOnD2XVN95VMZ+aIfQXbLi0gZsDHVq+MTo7z
gMoI8Kw01fErq8OBaYPHKCTYb+tZ3g1PXzsRDGNawqltHSTLpes4HhzMSie4S5GKQqsVwjWuOvaGRCw0ZwaQR+PTx8hFBvRrvQrHgS9TqucqW4bqUTa+VP4OQFuBO09O
BM+zh+zUAfEtGxg+YznVe9RYh0NXWNOmxk3f3J1dKjz5MWe6jrZ7Nf960ThBL9vrnoUb7dhzqzjRL9LdgvFPe/mE0/THssovMK3o/4oSz9nFi5iCRQI1fX9c8gM7hiRG
F4Ahl/oU2TgmWVVH5qJXG+PTx8hFBvRrvQrHgS9TqueA2YGB9KWjtS7NVB1luGVs5yIM9OdllrMKvacu7WJvC+FzcmBY5eLreHNcckBJcsCxGmAypUCUmakhbceNbK+j
hgH/dAW8KVhunehJ/Ob0aSTYb+tZ3g1PXzsRDGNawqltHSTLpes4HhzMSie4S5GKIIvfuN+HNGAtwCK5jDPpFAd4oahuQ0XIgJAeN2vQQ8NwcbsBar0WXgAUg0fzslik
U6bgO2hzpVM70iDAxRsbW8DI4k6l/Kxkpzgccw97EH9ep+M82DwKus07NE5gmiQYxiKaX6SGaW30rWSdbcZGnyTYb+tZ3g1PXzsRDGNawqltHSTLpes4HhzMSie4S5GK
ONwh3KSXuRoJ8ccbSichdtwPhqkfY5TiS8mNRmcslqLZm+SFe++dOD9F5YY4vA/L5yIM9OdllrMKvacu7WJvC+FzcmBY5eLreHNcckBJcsAAl92LLGRo+8bYEwTxZFsm
wSVzP3ZG0/U5OteFMm4UQ/ozkZVUU9VZw+GahYf2a3GflRzLSCGPe+MFhyieR2uf2qkkB9K8yVpiUp0dySzRfG5p/fmGqi5f9yuET/1k5KlI9nB+G0/kHbVHiMW/lsDi
lHSPOKfCKum6DWtcHWHfj2Li9wGPRgb74m0oe2iL4IUntD3HNc3FB8IeB1EtCQDmSw34GBtuCUygYGL+g9jmhZ9h//6nDo/tZePB9Sck7QDOKiJaDXqYCm6qPeSA53BS
bCpE4NSEBeKdgFI793ET0dSucPkihVI49lPNRtDRipzHhFaJK4XMe/BzInffZJoDDW3iry758mTmz8eX70BaiBwfA9Aq3oYN6hCnLT1VtOAf04hQsEpsAdId+v84GpAA
dnvicU+JREHfFXUywEeZfFW1RSytyEkPvyW9FRZctC4KPgMnB3rUqsbH3mMl9exaclkQjNT3KrFF+Sq5aKmiKDFdw0l5g/c0hKSKUhxI/Hmc4narxzYqqc7mkZCId4Ma
CwP8cCt0tnGfgFyUSzWhimqXq9LC5C9PVNwvGzDntSbwY2CTKtYtQzC9wwECag1mQujwxoUyJW7eHw04zF2SSKbnXB59uZ6zrB40jnkhwHh+fbmWDZ8TwYHFDZgDDlii
pMyqgotl9U8jhvjpyarO5wVJc3GXSmW4sNqC6VPni4mn0B8frYOh/s8yqICKHyselgoienRkm5V3Iv+4KYveRFTrWVl/PNTQh0C8h1JqC4OP+4PdXOzJjNw7XMUxMNDe
28EoxTkf4s3DwUrYpICQv54DGZze5w/y1A9WDiFQajTUJy66FSKqpKkQn5j2fqnSq0GAk0bmRG5bBguW1kV+EX3hdguXV1K8pU0dle17DvSPDWkNZ4dAagFDdMJdJM8K
VbVFLK3ISQ+/Jb0VFly0LmVjAiidGbO1KIIp7sTJRm7SViSfxBSbRFo236IEAIPnQ8wYiMQYLpDIv/lkzfo9CtMRz8Y5Qm5E8uVDfiEPmx6B7L8NV0FZGQaLjeQT+jb6
1l7p3HfM5qB/wCiCCDb5QantfaFPPtoDoyvfUjaxWi357s8r5xEUKs/3wJm8A1Q0rnYRjoLVcpr8PzTqTgvoVmx3dhL+bqKxcqOd5qz+B53FXeSGmDWkt2iWwF/WSGNj
0xHPxjlCbkTy5UN+IQ+bHm8RwvCyn2ub+KvoPSK7DxjUrnD5IoVSOPZTzUbQ0Yqcx4RWiSuFzHvwcyJ332SaAw1t4q8u+fJk5s/Hl+9AWoisdUM6c6cgSEeBCJVNokA0
Sw34GBtuCUygYGL+g9jmhSIJiFjmOsdHFaTrKeVR5EMNbeKvLvnyZObPx5fvQFqIB7PMO0kfYNx3qbXN3bVsEKfQHx+tg6H+zzKogIofKx57xPbAtO5vbhvCDNPwKtkE
Njs1j1W0KnL4BhjoV6t8mJwbKKF426zCJfwqh2QcaixWzSzRDm/Nw/lRmX28NtY8knUvHwj7pzR4PeUv7UTQgTFdw0l5g/c0hKSKUhxI/Hl/4aaKhKCs2VK5o9wAbS0w
aXunWyxHa9f0dU7mQdl0clUh59ERS610z74PKFcPQipJEuS5n6mHoR7nRNANTxViWUScgRhwWnalPNED5rxr3jFdw0l5g/c0hKSKUhxI/Hl/4aaKhKCs2VK5o9wAbS0w
ehKKNyN8Ofk/e5pBXc0QeFOm4Dtoc6VTO9IgwMUbG1sciyTPZtfoWaRw1Rj7bTLnAwYkvmxU+ApwMQyBGB8sFCTYb+tZ3g1PXzsRDGNawqltHSTLpes4HhzMSie4S5GK
5I3oEJwicf5mk85yCVZHyeciDPTnZZazCr2nLu1ibwuU0P3iW8LXiBe7mV4q89syxoUQWxdeVhcMqTG15aBrtPmE0/THssovMK3o/4oSz9nFi5iCRQI1fX9c8gM7hiRG
iIbGZKJFkqm0+DKyJ6qjewTPs4fs1AHxLRsYPmM51Xup959R91acVIagvumIbPMjTMLSu6x4Ia91J7WGRKayvAyEbC4nQRjazlycDJdkGHfATnCkUjaz3KNWBeacD8Ff
wdgg8VZlrm7gqWruru/B26NYKrHYbfWXtMRODobinFuajzMUHyRxpRKp9qkXVASVe9AJAQ9jLMccIDbyryxWWwyEbC4nQRjazlycDJdkGHfATnCkUjaz3KNWBeacD8Ff
awfUnSrT+sI22icKBRUnwqNYKrHYbfWXtMRODobinFuajzMUHyRxpRKp9qkXVASVO+P6KXuzmKQu5vTRlIHqWQyEbC4nQRjazlycDJdkGHfATnCkUjaz3KNWBeacD8Ff
DyWeJfRqXXnulDTl992mNUE6zXySCCMo3UqSg5Bp6a+OEfMyYXt5HPmQF3upyAS21kSHWwp7wbu/6JsZXxGqb4BKbTyTlINjKpIOR3+ZBvgZsBzsCe08DFD2k7h1QAla
jhHzMmF7eRz5kBd7qcgEttZEh1sKe8G7v+ibGV8Rqm+CUlyE5nVJzlzVTdxya90lwApdfrcKTv6PuTHpfHsrHXiEc10TSBM0L49fGs0zdFI/z4wSe+MrLDH4lwJU6A3g
7CPnEMXAYIKurkd7BZfgAUMN4PSPcUN5UaU3Wq2lq1ryJGO+rSjRl3AeuzqsNGyFWBhZoh7T3oDRpfZNav4SXgTPs4fs1AHxLRsYPmM51XtHtWffV/a/nQDDLRn5KJOU
xiqdcNQeFJfbQI5pO5FX7NqpJAfSvMlaYlKdHcks0XyG0j9W7wwlpjCqFvhZkCwU0m4Ko+tR/ylwXuNI1qHPsaIEmdbCgMA3WLbPZTcjvx1ErqrRWguLLMviEzmaZhjH
mYtJ4KB8mZWY+vKHNLPrqyg+vrW9xFhmrvHetGFVZI7HhFaJK4XMe/BzInffZJoDU6bgO2hzpVM70iDAxRsbW8DI4k6l/Kxkpzgccw97EH8yl25WTw5UKkKPGn/CWRIW
GL8YNP3qOXXSIB4Rj+Nj7r+VCzpbfEAaFX7dYj9tmGY6TnrhdQHpMIOPU/Sy6mE7c8zoOFdJccteiSMYYAhtBlUh59ERS610z74PKFcPQiofOq4ypG/J4ISgKU14U3kM
IQc8jApCQTq2VAro4STaWrhPVVSc2IDdMCgX1Qr0T0jdKpH0i4bH8uAJY/pXzfjJF637nXWg/DhjAeLtTqzIAU89XDTvBbWdpXyOYk7GaNH5hNP0x7LKLzCt6P+KEs/Z
xYuYgkUCNX1/XPIDO4YkRpGFiua4YOBfOEaesosIVlsCjCUa+ijpbYOIRgSqq0owhtI/Vu8MJaYwqhb4WZAsFNJuCqPrUf8pcF7jSNahz7F+tXdFKQCVv+PSoJRmeCcY
chTn6sdGyr1l03TafB50SvnuzyvnERQqz/fAmbwDVDSb6gALVAONht4MM3eY6e3Z1K5w+SKFUjj2U81G0NGKnLPR3uURSNWzbzcV8PIfbtrUJy66FSKqpKkQn5j2fqnS
K2IT+xbUpmVp5mrDdgq/xksN+BgbbglMoGBi/oPY5oX+BhttWkmBfN7VfNrTUF4tNjs1j1W0KnL4BhjoV6t8mOz7lORMOdyNJiNX7mlZbIOPnz/ngp7PKjRTjQ6Pmbkh
JdtB1X9J8kGeQsOHFgqxWjY7NY9VtCpy+AYY6FerfJis8gCTlEBT/A2lMJw9b4Lm7mTC0TZp1MlFWYKsyN+7oQ4uF/QV0FCXC9KFVdHfV5OkzKqCi2X1TyOG+OnJqs7n
ju9a/ozOKvEV1DVUpcONorCiXw4kZajYIqb6+Nno6+vWHu9Ft5iS8fbD/w8RDqWWMV3DSXmD9zSEpIpSHEj8eZzidqvHNiqpzuaRkIh3gxqMAIcXFww0l91w10fxDQOq
xAL8OW2A2ssdEOVVHJKOeL7vwP6ZfuUclAiGvjTCURWNIPcK1p+fDReap/Rig6guVOtZWX881NCHQLyHUmoLgwQjD7xPNwLWgC7FNrzQj/yMAIcXFww0l91w10fxDQOq
xAL8OW2A2ssdEOVVHJKOeL7vwP6ZfuUclAiGvjTCURWNIPcK1p+fDReap/Rig6guVOtZWX881NCHQLyHUmoLg8RWrM+ky3ptwzZCKQy5wK2nrnQ67YLWQiWFzXCRPbbW
0SihhurbG49Zar8th2tD89QnLroVIqqkqRCfmPZ+qdIutlqSe00HBtFqcJAeka9DNYaPlTl6KnlYGLsn2mcq6Q9PcGWx9IlRTapZfydcmNqLMfp4XzHaFGLrIu9nDg6t
1CcuuhUiqqSpEJ+Y9n6p0hc8OYXhL3jVrmI1RIZkQ5li4vcBj0YG++JtKHtoi+CF3mqf1mKaEIjwnLFVsGZqBb4oXyRk9o58++Qc9TdHt/gmmm3ITT5Sri6eVw107DdN
9qWo34TE6jUgmnBojggTbqTMqoKLZfVPI4b46cmqzueO71r+jM4q8RXUNVSlw42i8sPN4SVPWxL2wHsa9KUpBAO4Ao+PMbQHFUN4kXwX+NuO71r+jM4q8RXUNVSlw42i
akDHEeQX41wb7u2KHtUlBs4qIloNepgKbqo95IDncFIn9zAMs3c5wgPj8Xv+o7jWirQNMUnE7I9sXrvePZ2Oio7vWv6MzirxFdQ1VKXDjaKake2Lave97O7oz3O5Sean
Mf+yHUzi9I7nY1ppt56SNtMRz8Y5Qm5E8uVDfiEPmx5bBTyKWPBgoJHwuxySQf3Bj0g6wXfJCamY3mtJjJdxE84qIloNepgKbqo95IDncFI8Jbj824BNxJX9x0IQllwk
2qkkB9K8yVpiUp0dySzRfEGXy/STrSZIASilcZJPswJGoe1KvKTR9mQfWH4cWj9AiPIEdmLskGlHVILtPhy+lc4qIloNepgKbqo95IDncFIsKXIC+H7Bc4RIMtzUZEts
KBlUqqzcTtqU4zqDjAVqDwicC98iNqFyFhP7zaL+Qbe/JU1TlhyqIfkss6ojS5Duy+1lqcSxIu7S8TwdbRHWSkSuqtFaC4ssy+ITOZpmGMcJ8imp3qNzXT8cupIVdfwP
OQbfwgq5cuxNbnGvNgMlrmRcNwQ7ub5FuxILF2M1GMq/RVcMyqT+aeKzfmzaDeYCt5kkny0gEXKGm2zCIziQ3/Tog9oxpNFXaMiVstlPkjIxDmxUNcQqTZnaBbLti4p/
okiZvM70sM1kay/8QwD8u7Q9HHporetd0gibXCGUn8brCeZPVj0lQ2NO1kCKp2XPSW9NF6CKBuHLdrfZ8dEq9qQgLfaVW9wip5l5kSqsCgnOMywmofQzuM5YrRxCFA22
SBlbEq0KK9rZyP8kp2bGtmRCrLYr1iNl4IfUMQ/Yqv4YGKFUHp7gGOm6D0t0MQAUltBThPnJ5gHhVExYuCzcLmRcNwQ7ub5FuxILF2M1GMq/RVcMyqT+aeKzfmzaDeYC
d86BHbgYYy26cK8GFILP+VOm4Dtoc6VTO9IgwMUbG1s9lB4UT+TrgFLlM/SYQubAOLbPO27P/Isc/D0hcQASBCTYb+tZ3g1PXzsRDGNawqlkQqy2K9YjZeCH1DEP2Kr+
GBihVB6e4Bjpug9LdDEAFDu+ktBT9WPZjkQhjd9LeBffygSDugamsneJinKBrcqO24c+3UDaZ2oNEgZhHQgzHvu77M0VLOcWoWKpxJ3O2nZvGziWlZ8ZgKsoSwKoiJfU
KUQ4MOY8TOL4inlOOB2rQ/SSgYmgSh+5ss2Q5xP4yzHLN7YX8UuyWKhMcjJkSR5ISW9NF6CKBuHLdrfZ8dEq9uYWHLpOtY+VwYepZNdfUd4WJGBqKabhfiSYdmcS35ND
I/yQCMF12La430Nk5Q8acSlEODDmPEzi+Ip5Tjgdq0P0koGJoEofubLNkOcT+MsxqGnxrGEqrxw/rNqfPkHAv5OMTCmJXv4mxAD6f2auv80pRDgw5jxM4viKeU44HatD
9JKBiaBKH7myzZDnE/jLMWDGLRE062LN4jU4RDHojBodN4eMaXHZiTDJNFsUhGsXrizvr5OTPRaSaxKTOXKv8dtgQeVRbawt2RtNh3iMMdfyNekr8UBA196vItGtVJ+j
GbAc7AntPAxQ9pO4dUAJWtaPD5cDIrRUHT9uMwCaPT8MBF4R0XjuPq/WQPKOD54GBVWqzecYaqgKQLPJqwVesRi/GDT96jl10iAeEY/jY+5/4U25pCQPg56TFSw8iK10
81gbO/9sMm1VAmmPp6+i9DPA8V240OKQrUZ6YFBEEWkk2G/rWd4NT187EQxjWsKpZEKstivWI2Xgh9QxD9iq/hgYoVQenuAY6boPS3QxABRrgUINEKEOSv2KGQCvtp/4
RK6q0VoLiyzL4hM5mmYYxwnyKaneo3NdPxy6khV1/A+y4aBji6WrZpfZgoMszWEjN7PCaLI4cRjhIL3vgwtecvmE0/THssovMK3o/4oSz9muLO+vk5M9FpJrEpM5cq/x
22BB5VFtrC3ZG02HeIwx1+EdOkPNuoVLkGmaxYEi1w5ErqrRWguLLMviEzmaZhjHCfIpqd6jc10/HLqSFXX8D7LhoGOLpatml9mCgyzNYSNzlPRvzi9H0JyWFdePQ63k
p94Is0D3DznXE0voEzpiiVDTCdO/GdTQopNwPNAhheBkXDcEO7m+RbsSCxdjNRjKv0VXDMqk/mnis35s2g3mAmYmYB0z5dqydqI27Fe0vvXdG33T2WTp3w6Xufevs7+i
T79jZcbf97PBlsoX4ec8sfYdO3i80/A9VbIA80mdrM/DThk0HSbbuy/SuJkQkbxpE9KRpBPg/w312VdQqPuQwVGHwkJPoaMWvnxZ4Z4/0duLrwScwfHp0KyMh6BG93ON
GL8YNP3qOXXSIB4Rj+Nj7n/hTbmkJA+DnpMVLDyIrXTzWBs7/2wybVUCaY+nr6L0PRWk3ypG+O4XPSqdKxFKtqrM/YV3Dv0o+K/aninPxDDz3TrBj6aTgkU7z6wtygHA
KUQ4MOY8TOL4inlOOB2rQ/SSgYmgSh+5ss2Q5xP4yzH4vqbaex1xMqd2JrFuHvGaMygrJvYQ0cwgt+9Atl8oZOE49NW1ZCJkp1K/wLyRxJyMNovj+eSHfwz5jOOw7FLH
YQVG1ckMH841JaIiS9iqZQLRabjTqKKEkhkdWGIZOTFSOli3BozeylZcYh7as8iRgitDv+xGxhazy7VMRp+Ufq/PeRY9Hmg4JV/y4PqF59OQjUaAS6lf0uphZ711XmqX
TH9cEBbAs58BcWz6FmT06iHp8VHjQDyNCMDGQXhaTrzH07rfLPFdbYNvtOnqI+K9zqFPgqjAhTJs0Yv4R3l4x8xjBsAeDwX2bV3QmbMB5nY3m1CrQlrwNJbBsjUSjKNE
NvyK4lRdgFV5R1kYyNE1sXGS4V/vvvWP2Zcvw/q7k0n4VvQA5EzrI3+XxAK0MHupJYNkUgkny/BB8vutG++PGzbpS9X17fM87rB2yFxdk7YCPFNnWC6EuYklRjusNcP8
EKrfL5rI2smvXWEy/ZZ/zF2vtErrds0n2rcZLeaVw9TsO+1gbZQCwPzsUo8rfF77cZLhX+++9Y/Zly/D+ruTSUo+5LeoIlWPikeanWDIPttPRqPk4dvo8CgRcVLX9Jp3
jTL5QX7edooZR1b+QrblcXFHx2DITliQ8qwqaYxZsmz8suPq/rJ2H+Qps+5c1qUWJUqIi+oA3Sb0lnxVsw2q0iiWFdiGatMNf/DSy4Eo8XwJcTpJAzODub0ge97tUcEE
91H6Ru7CN2bq9Mij/m3xWD6X1GVjyasG9PGZYLL59oT2vgaL5jBjzCOTpPfXupAFzPe0rVq2Y8wJ+KauqKmpSab9BjJ6gDZ79bYz2fDAckglaHVSU8T2QEtZzfYTQnca
w1Et2bilAA0I1UyxtUVyYxT16ChVOYHS0+kRPH+caY9uFWmvnd1zPwYmDu8h4vA3CXE6SQMzg7m9IHve7VHBBPdR+kbuwjdm6vTIo/5t8Vh4tcFphT0Ip50YYDdSdfS+
VNAJClwEzSRIQ/+rj5l7TKHn42T+XmJxhnBRTJhhQef2vgaL5jBjzCOTpPfXupAFzPe0rVq2Y8wJ+KauqKmpSZb9haDSWjJn3x0fHJjKR5xyBlWB7McnB0qm12ec+RFR
C8q0oUZ708uamuqEe9Xb16foNM+AKWWS57NiWBoHGJiCklAfLwQ33Z8Y+j/f3xcRSLyAXtxA5A9ADJ7RIKI0RAhUrbW8nMZohwi3b58nrEudWHTroDkxeFmyXUX5fqjE
9r4Gi+YwY8wjk6T317qQBcz3tK1atmPMCfimrqipqUlpL2u7n7SpafSRAkrZC8oJxhDfM/XBc41ox0HUlUVAkkhQ43V/Eziz61QBeKEwk3ifKgttNbycqsmJug+Yw9wG
C8q0oUZ708uamuqEe9Xb10c7x0tl9fVclK7QOaT1Jb5xiWLm+5xAimvAohv0XV52FPXoKFU5gdLT6RE8f5xpj10WeRNSj2FtvT0ZtfwTFFtNGTnP2o/O1xPD9eBsU3Z9
J3Fpnc3sxC/tiplq1keawRp3pdjhqocLZduAP7gv+QG0LpPfWAn2w7CdlUvbrdskUnJINKOYscfcdAK3tP14XAvKtKFGe9PLmprqhHvV29cYA2Zvq6O9jHO5ct9d8cJe
i/aUZ23UJYsL0c5qEHtf2y2KUpGiqla3dh7es4K6FiubTTEoTSdfPX9A7sLJ3flAFPXoKFU5gdLT6RE8f5xpj3u80LLLS6sADDh5RxlDYZyddZa5nnDBA+tIErMEN7bA
XtgJb7lTTNahwPR/5wLlzU5oqtolIpnAiX79xJOAO7bEOFNSKmsHDs9q6zOiUBb8SQhlP3A/mQaLAue2+2g+KiZsXNdBSKzWMTuTUGQRPLR2bxpHfjTSVHLRf3I6cSxo
egAKMkhtg3tcDKmldlg0mxT16ChVOYHS0+kRPH+caY//+T8RAoGc/pPoElIoUxnu9Z9siPY85FEKuAMbW0MW3kXGLoSgA/CfSmQ7HFWtGmrn/kmKZ50eTcwgJjqT0/v/
XtgJb7lTTNahwPR/5wLlzU5oqtolIpnAiX79xJOAO7aWOf1XSWs0gqj+uzI4xkBAKxTOl6G+1z2Q5b2R5Dh3XOK33+mitoBdTqqU25mscsiGVVw6AtzjF7asqV7YOS0J
ta/D6gPxv8DM9iITA5t75Gu3gAS+JcWajCR5ccmQO1tFp0jpoBCR7RTLpXWhCuf9IbQFRN1/e2u+ra/MyyXHPl7YCW+5U0zWocD0f+cC5c1OaKraJSKZwIl+/cSTgDu2
EBZnBV7HjFuOa58Lqwhy93Og/FnN0keH7XeoY36L9JixQG5nbk/pVJqNEWzS2t2CCXE6SQMzg7m9IHve7VHBBPdR+kbuwjdm6vTIo/5t8ViRI2O2OVIlBuyjkCExhLkh
9r4Gi+YwY8wjk6T317qQBcz3tK1atmPMCfimrqipqUlPo9ummtmxJHCnEnUnurg/aAWYcouPOKYIPXcgrHVuR/rLdwKb2+HpF8LOofMZRZS7sKqk9Jw473xs6bc6xc+L
TEpvSSWvZEO4+4UrUaZf2shJVb59+687ImoOFPgUIA52bxpHfjTSVHLRf3I6cSxoRBk9r5Xx8tXd9N7Lwd7lkSachb819HonWrt0x7GXbk4yK9FnJF0DC/WZOnoUjH34
RlcCtM0JBeI9iwY5Cz1fCQOo6QMjK/tEfF/H/nOuznqDFQYMhM3IB7xdZw6G+EoHUSMfBy7ZnQmWiuD1URK/AYvTfrTLSqst0XcFv2JHOd5T3f7LXYSLfqJUfneAXD62
IxJxePMmsVH0/u9kp4bxNvBOnTOZVyYBJ4Td6KWF+vB+hs7iqZFrNZ1gxVNZcV95zPe0rVq2Y8wJ+KauqKmpSR7K7eywiinHF//ToqRZK6uL0360y0qrLdF3Bb9iRzne
U93+y12Ei36iVH53gFw+tlIR09NXh/Ntb/qx+m1jaRYiKf3/kOU3y4Lpu8E7BO0onvu3guyz5dX0h8l6jEW18isUzpehvtc9kOW9keQ4d1zit9/poraAXU6qlNuZrHLI
63EXfUZzeY3INQ6aCuUDO/cwRJFEMb83DAiPYzYDMspqxp7RKs8+ohSU18s0XEzAwOOWDlCNn9lmc/4xMrqd2Ny93f8X9NoUmYewWHADAkpOS9uMQKrId/FHvU3RUZ9H
i9N+tMtKqy3RdwW/Ykc53iIXBGQI1Av5wcSJMMoh7P/ISVW+ffuvOyJqDhT4FCAOdm8aR3400lRy0X9yOnEsaPio/l8uQKbAhEVZ+0MJHlSwaHVWPBl2nPo2gVCFWTNW
MivRZyRdAwv1mTp6FIx9+EZXArTNCQXiPYsGOQs9XwkDqOkDIyv7RHxfx/5zrs561l4ftzd3ff7k64FiFPDBs53XpfnqudT5m1Y0ravV1R2L0360y0qrLdF3Bb9iRzne
U93+y12Ei36iVH53gFw+tpBR196z/rpWOxUoqS+Oi8e5KTiMRBIT8+2cQEeabdwhfobO4qmRazWdYMVTWXFfecz3tK1atmPMCfimrqipqUluxqiXj5WwJ4HmEz7KSV9r
i9N+tMtKqy3RdwW/Ykc53lPd/stdhIt+olR+d4BcPrav1DF5w7r9xK758KYBmR2HwEjJzQ+vguoJ7aIBfESGAp77t4Lss+XV9IfJeoxFtfIrFM6Xob7XPZDlvZHkOHdc
4rff6aK2gF1OqpTbmaxyyKianILjR4fXaQpCOFbwKi/2vgaL5jBjzCOTpPfXupAFzPe0rVq2Y8wJ+KauqKmpSWLbVAizAaOTO1ANVNEINXFmD6N4mAK0TdaGgrCa1csk
+st3Apvb4ekXws6h8xlFlLuwqqT0nDjvfGzptzrFz4vt6MizDiZFtiRdF87dAeCwGLhvwD3/bS5gZxDjIJrNnWYAOrcfFNRG1LgzLoh87x4UkwODos8DMLaLaltLeYNu
KmVT9sKa34gzyLzGOCV+gduH6Xy+I9nj5NYBsnGG5HrDQxKuAc1PhEqZ6KJdPpI1jriEUaKCbNLG/fe/9dtJlWbH8hrx6zgiNBmacZZ48akMhGwuJ0EY2s5cnAyXZBh3
48KjfcMSwRHh+h6stVop+5rNY96LxDxbKknZohg0rE9ZOGFKjEONg3Js24m1eZiQVjo/kA2REOsbp41a2hVhe1Om4Dtoc6VTO9IgwMUbG1tyOFg3twEndwyGF3UHcrL+
h2qx5VEoacGAOMTyIZVsSoN+WhtAr8rjv5FiExR7CIyJRCUYAHThVdu53iUlDy+05yIM9OdllrMKvacu7WJvC14UNKgws34GJsVaRV/+mJG+8mm5Xg3iJoeJVwvkrQ3l
caxCVjjDXntsopWrO2r2lmzVFar75CagUuaDiSXJzg7fqvrvXqgR0nE9VotiNodQ/pSHMoFnljdB86Srl3rzZT1s9z9bOO2+RusNsQ0FoXzCy/YI7g/sZZuvuyKzcLX+
WThhSoxDjYNybNuJtXmYkMvCUc90x1uyyIqzT3Pxc1YZsBzsCe08DFD2k7h1QAla8PUZrvwHxt2PNViA2nWv2p4WQMHKYRFCuKeggrJC9+Kzj5q4oOkNFpoCUPCWc2hi
PWgbOdHuPiO/JvGQ7xmxPyP8kAjBddi2uN9DZOUPGnFTBmoWuZy0yJa+iGXEQZ9FzqIXJujmJvgUvwTFmUbrJDZDEASYRD9NbEgYG6JmCtwWS0YhXvzxFa+RjJNBpr8J
VSHn0RFLrXTPvg8oVw9CKlwUhfnWfwsEH1cfttm1iMd06fBKpSrDN7Oo2evx4BTjKLGnfCxH+7oQpbI2uOZJKWRxuJQDwu8AKgL+RpHzfqxJb00XoIoG4ct2t9nx0Sr2
5RDNYnF21wmtKyV0txEhcc8oxwxhq9Ib5mKIG72IP9uAO8DMVmmlsgk3CiXAdgnFbjLu7TrHPnOpS+uSZGdaqYv+z/HuxEsny8q6WG6duGLyBmOK1Fw5JlexFny+Etez
yC1mUKaFoAN9o6/R6AbxYuxwKPn8Hn3Tl0SQX1cEUnsacI4H8AGy1hg88xVJFsR+FvC/cys0N2Xi3jAPUpwFCktoybDiruuML52iuyAaIJtV2aDBLZgTs/r5rAXOydpv
q7d1QEie7SBBS+S4/YLoUS+iKXD+XZWWUvS1DNfxdXWf57V5hGbPEjYgFY+1AuvmMr0Nc9JW4GB9aNApi3IGi0j2cH4bT+QdtUeIxb+WwOJv2w/Tn/Lcb4Ae0thTMKLP
P8+MEnvjKywx+JcCVOgN4KDIJNMbAyBfnYlMnAMmCeI2ipEDfaPplA2ubiTbB831+e7PK+cRFCrP98CZvANUNAYujrXVlhqtpmMgy1jV6kDhwMTkJg97z7Px2psnSPF8
+e7PK+cRFCrP98CZvANUNAYujrXVlhqtpmMgy1jV6kBIcLaoCufbryO+23p6YkCBVKpm/ZiI+5Lm9ngKVSbcMiigy/VvIf6lsU0CZ0Ua1dXOKiJaDXqYCm6qPeSA53BS
Fn9Y+zmDdADkdxqY+j+MrNW7H3qS9Kbi1CG3u2zgDZaxeB1aYBEhpzFZBeNRLDHJMV3DSXmD9zSEpIpSHEj8eQ2AUbE+EFMeiYElkfqezYjk2N5yF5jck+yKgcorncTr
U9V0sIqRrt7JY2lKiAdYFAO4Ao+PMbQHFUN4kXwX+NuO71r+jM4q8RXUNVSlw42iuHbE1sH/1ejf9uC1RxaWCxThfDmh8jujomvjKAsvW8/OKiJaDXqYCm6qPeSA53BS
Fn9Y+zmDdADkdxqY+j+MrAqdnomrWSEteYRW7b0C/iYeFaTT3ZF7fa6nrgmI0227+e7PK+cRFCrP98CZvANUNAYujrXVlhqtpmMgy1jV6kCcRS3hQmOaBh1hWgdTMxEe
MV3DSXmD9zSEpIpSHEj8eQ2AUbE+EFMeiYElkfqezYjk2N5yF5jck+yKgcorncTrH/FPkCjRMDindezSxtC/ejjQaDY3Nb2Uv7DyJVsyXsib0YHuRV46oGHoqLpquHRb
L/f9MX3DkCmM5EhhqgGohdqpJAfSvMlaYlKdHcks0XxYGZyUowpZpFCWhtplQ6fcw24CNW2Kf3yAc/afDNoctBEyMmh5BjMlLRrMfgNF+Z82zZGmY/n1ZewiHH07BXup
h/kK/E3FHoRrytPcao/kh5Yp8R5iOx+/1c5KX06kevQ5Bt/CCrly7E1uca82AyWu8BS5uSJDI70Hf9wF9QmY6o9b7Cm4EP69t8NgWiaVPVRRYCN7DKpwzdbepFBE0XYK
tfbUomdAiazIfTTylvlK5zKtcQiJf1WZnZxtTmQnsiH4bOSSMQ2D0BjrXvKwHbwmOvl+g4CKcd2n20BRSs17u5iFkfc54PhfkfqEPX9E2BDDB6IZJykGnkgrRbXLc55J
ONBoNjc1vZS/sPIlWzJeyJvRge5FXjqgYeioumq4dFsJBYOiX5QBLQcd3I9rFrEOq2IAgAscY9wzlRIrTaBIrYie6h+l6j8oesWpcF7Zg67AXGeWmG8DVA5m6dL1HzeQ
JVKa5rWhGmJUyc4UEEuVCMGHyagQmT4BTo55E7qaHV7GFxb1WSsPzO91vpbaowNuE7a3/OLXwvOVe7KnRtcg1rIs5KFt9+9424bRKSSyUW836KnGGJOFNr4+G9DHFkX7
/YgiSz/i/Eu267YIlzljoMmHtMaA+RilsMAeNqM4HYYVF7wyx9on/eWFQRwzqlQJ+BwVw5/Kir/s14M7ZhJTff2IIks/4vxLtuu2CJc5Y6DJh7TGgPkYpbDAHjajOB2G
P5/o93WhNQRCFp5YUDTPr2MTxTelA3SLFuSpwqwevArfjTs6cr+bue+Y8trbk3YLi9SoZlarFqPNkOQaRqlMrvHtjdciwTsiagX01o0HKdkVE50PFNojPvIbjqhsPFZ2
/YgiSz/i/Eu267YIlzljoMmHtMaA+RilsMAeNqM4HYY/n+j3daE1BEIWnlhQNM+vHL6Vvz9bYjgmsGyvUT0B3/2IIks/4vxLtuu2CJc5Y6DJh7TGgPkYpbDAHjajOB2G
FRe8MsfaJ/3lhUEcM6pUCQRYKynxmQtcqYitO9SDe/DGFxb1WSsPzO91vpbaowNuE7a3/OLXwvOVe7KnRtcg1rIs5KFt9+9424bRKSSyUW+aMzIf89pa/PREZt9ZHTsj
ZMXH9z2JsBdAKGFZf/unYl8rFr5FDzyrDI2HBrzGMzWorXQ44JowOtnNk0KYdN3lzioiWg16mApuqj3kgOdwUkq7wSZ4ygLZ6y0cK1hbJPcqZIMkfLfoJGzgVoW8yiCb
6fFQUphumhz4jjMd69UWwpmnjUtzJWvZWN8tpdR4M+zfjTs6cr+bue+Y8trbk3YLi9SoZlarFqPNkOQaRqlMrvHtjdciwTsiagX01o0HKdl+0vUFIrJSPr1K1t1YhzaG
3Rt909lk6d8Ol7n3r7O/ovnuzyvnERQqz/fAmbwDVDSCmWghXUGKuTf1YfK+bWt5s8mr/fEWq/sDcTLebnm8Oof5CvxNxR6Ea8rT3GqP5IeWKfEeYjsfv9XOSl9OpHr0
suGgY4ulq2aX2YKDLM1hIzezwmiyOHEY4SC974MLXnKkzKqCi2X1TyOG+OnJqs7n6k/APdVU5xndX668+awTDYjyBHZi7JBpR1SC7T4cvpU40Gg2NzW9lL+w8iVbMl7I
m9GB7kVeOqBh6Ki6arh0WwkFg6JflAEtBx3cj2sWsQ67bs+NlNQF5CvKlWMj+5YdFPLAnekLoRSQ0rT9BchzEdQnLroVIqqkqRCfmPZ+qdJrfvN+FjRq5ne4TfmmTdBG
boxLiFr4gmWaiTa3aWnz8yi9Fuy+czzBxFxoBQicMYRp/fSny7c/o+nsT9GO8iHoeeCmxIetF3RIro9e9fBehKRyuzYkNY+meLV2HUienHBU61lZfzzU0IdAvIdSaguD
qNGp79sCzjbsLnJ7HBgWq+oDBb4wwct4yOXtGYqHNbWRkWVmaXx1uo/fNh68H2wfvGGmSNB4ezjwyuxCN1RxLSjuKOktBsg797cFGUDA0EDMBYWMoAABjKnD4bRJKNSy
cye8RBdQ0jmK1lSuBgqUprm8K7/j3kuyyjIkWCT6hWZiXwSqpNOfH4lj8DuGxmQQZhaM/z2ptoPOVzrMe+tO6+g5HWuKxsdPKfwQ0G1hNNr4ybU8+t560PoQfj7ofU1R
MV3DSXmD9zSEpIpSHEj8eXg8vH86wRFoFp13gcXAMbVwXQbysSkuwBD34KILrmMlzioiWg16mApuqj3kgOdwUsrVuQn5gAef1we6gAmcvyYU4Xw5ofI7o6Jr4ygLL1vP
ERUGIDzjAGNHZR4Gh8drqgIQX+fUyPrGDjdEabLla9U8GZHeeBf22E26p8rR2elzAlVP8gK460g8fqvzg9zNPVUh59ERS610z74PKFcPQirZsU53g3rYeb9OpzJfxqrO
HKlue9FFcRkdMJ5QZh8JwG0dJMul6zgeHMxKJ7hLkYr7DdNTBouIDyd+0h5pIKvKtx4zuVyUbBtjI7D2ID5rKSTYb+tZ3g1PXzsRDGNawqmOuIRRooJs0sb997/120mV
3n5YpPJuvtoHBTMiDhW6BkgZWxKtCiva2cj/JKdmxraOuIRRooJs0sb997/120mVqL8AB8hGSbY8AfiBFcQfCUlvTRegigbhy3a32fHRKvbOEWM5qgin9XeKcW6V3Scq
wbNxf8cbsI/cKRUVxOss4/mE0/THssovMK3o/4oSz9lse+BqCcjvVxI5s++8i7jhCx4DrqhyBfIgOQf7CEI7T0lvTRegigbhy3a32fHRKvbOEWM5qgin9XeKcW6V3Scq
wbNxf8cbsI/cKRUVxOss4/mE0/THssovMK3o/4oSz9lse+BqCcjvVxI5s++8i7jhEb2eKKa7rHpcdW8cPNADnFyjdgFlFjzcCggeor6FXyj+lIcygWeWN0HzpKuXevNl
AscK1qwacUNjy9iaqL7kaEZIm3QSM+vAVLo+JUPzj9n+lIcygWeWN0HzpKuXevNlAscK1qwacUNjy9iaqL7kaHl/FErg/qaryrI/HNwcPvVErqrRWguLLMviEzmaZhjH
UQwj6rQdNhLPeuPrtygcRDWrjtqdIYZygZYH1Vw7qxP+lIcygWeWN0HzpKuXevNlAscK1qwacUNjy9iaqL7kaOBZZijJ1EVXdjw9RC0V27JTpuA7aHOlUzvSIMDFGxtb
UQMZHCN/OoSrOGMyHyERrR2hSuHW5vB6RW07B3OKTO1TpuA7aHOlUzvSIMDFGxtbUQMZHCN/OoSrOGMyHyERrQGxXzsqJKhcTK9U5X90IbsNXX3VKn4jiMuwMXFr3QGf
Prdxmnc+peDSgbAz+JjQpEbGUtN4oFy4U91X+bKzI3qsOBxp7Ockz5a1S2udZx3cNJHWizosdrRLmHs4SjjTbWHmQc70JRIAWOSKIwnS4I2MAJT8317dmAfsqhLrn6Ft
C4pawS8VL4qX0Uao7xEfr2XzZSXzHNbq/yAGJlujqjejseuc3nJUjzsBaZRVKCITC4pawS8VL4qX0Uao7xEfr+pt5fYFgXGhC/j93uCfMHGQ3g43kPO+mi2d91wyXkLd
8PUZrvwHxt2PNViA2nWv2uSPmfnzPZQ1vvV3ToYs6NJVAtaRdzcVQ0ua8Z7B2BO4C4pawS8VL4qX0Uao7xEfr7yAJlbaCENd2xijg8aRizpDFtWXdNTVoXZvZ1++CQlA
i/7P8e7ESyfLyrpYbp24YnFeDkUN+0tzIKSDsxZ+QByW0FOE+cnmAeFUTFi4LNwui/7P8e7ESyfLyrpYbp24YnFeDkUN+0tzIKSDsxZ+QBzlopivdtYzksNqyiC8GXJa
5yIM9OdllrMKvacu7WJvCw4pvkXo6UofgKTU+T5Izvo1ho+VOXoqeVgYuyfaZyrpi/7P8e7ESyfLyrpYbp24YnFeDkUN+0tzIKSDsxZ+QBxX9IeODYn8/+62FSULa1OE
51n2OMQKAPKLC1iQO5tAi464hFGigmzSxv33v/XbSZUHNG/67ZZJi+WUBuZSWp+w2jhutWSg024jL5jPiV6cPFUh59ERS610z74PKFcPQiouccpQkrr8MiODFqt5gfrP
QLfcNwWVyqlTPFJKx6pcOaemElHCcrTqPp5HRIEna4xTpuA7aHOlUzvSIMDFGxtbUQMZHCN/OoSrOGMyHyERrcNOGTQdJtu7L9K4mRCRvGkux14n/JoC+KSbEH25dbYe
1I7avMtgryDQY3vGHp32rKDUVFFDLvzfNOrQvn5Tnfd3fxX8o2BRfh4M86HnCqb1GbAc7AntPAxQ9pO4dUAJWvD1Ga78B8bdjzVYgNp1r9pG7QpbGrHlZyHW4Pr9oGGW
asicAL8gqJuuJfJ0Ds2TdOciDPTnZZazCr2nLu1ibwsV67Erw3SrSlPBiRzUOl8uqKQ7xdDwFvvyXN54OdlDy1tLP3b+jn0N8RZAPZ0QV6BVIefREUutdM++DyhXD0Iq
LnHKUJK6/DIjgxareYH6z0C33DcFlcqpUzxSSseqXDneyJCdg40YLR8y0th2HuBqjriEUaKCbNLG/fe/9dtJlQc0b/rtlkmL5ZQG5lJan7BtMMuN226dJ/btcAQiufha
GbAc7AntPAxQ9pO4dUAJWvD1Ga78B8bdjzVYgNp1r9pG7QpbGrHlZyHW4Pr9oGGW3BvvA7rZr4725zDhsk2qjuciDPTnZZazCr2nLu1ibwsV67Erw3SrSlPBiRzUOl8u
qKQ7xdDwFvvyXN54OdlDywdDEYkMwnRvk3kaLX2KksdVIefREUutdM++DyhXD0IqLnHKUJK6/DIjgxareYH6z0C33DcFlcqpUzxSSseqXDlXI+YzzVdyxTbobH73FBwF
1I7avMtgryDQY3vGHp32rKDUVFFDLvzfNOrQvn5TnffHIs9UhdICX7rz+RK5pG+aOHWYt24mOLqMQVGMeiuatMAKXX63Ck7+j7kx6Xx7Kx0RMkcAK2W4Q5W4NFE2gNJ0
gEeb8SDsFbkp+aeRR/Q2uGx74GoJyO9XEjmz77yLuOG32jVw8+q6jSyf0GXvz2a50RUIZUx4cx/SBc+W3ZK/QgyEbC4nQRjazlycDJdkGHc+t3Gadz6l4NKBsDP4mNCk
OphwATLtaA5C0EoIoK1V9H3cqvH/E/vBCCBSsn3I5qBDDeD0j3FDeVGlN1qtpata/7rQJe5DmFW8F7GMekyNfmzGDWfnIrk/ihyQtyyn3dtS5fMeUwGSJDGKBhVmOymU
2GkGfN6uQep2GS42KIyHFvowe4jnd8hxZKsqYPtJ5/sCkImqeM1C2hN3uzTxjhC5fO7xLf+Uu/HMZiqoJ8Q8lQLqHGXEYhCfbIHG7y1d2rZtZFLAXPmPCyN1DhQKjFH4
O4G/5U9ouFUo74mxTU0PiV1e7eD6Pm8aAbsqeBO+NYXjLmZY4nVyxw7Q2/mMaCw4wGQ+SY+m9jzCzCpIMm6XmbDc87kTQZ7FyblToG6DvJoNnK+6Ck+YonyygX7Epq74
kzLpU7DtH9Ma9rCM4EUUWgC8cDWNyr8LBgQCgcnRe4ExsUfkMkvKO8mmX6YN8HXiBobYEQ+Nh06EWNOfSwHiY942mg+m0arPzU1+xuuKP4EFK04fBmDzH2IzsziJx60F
ys5+d1LWLIUzk8A4UjJClD6e9H2nLCrkZgK8gQzlyNA5+XSKCIVHX0Ept9/xfcre/tE9iETXEsQ4MXKK9qKVhrRfr8T9oNdZ9sFlfi3WegtzlRF0lz1AduefuWJ+p7Pd
gLpbGlOEEtOLDtevsnT+krgMg4osYXaXp3d8iceq2t9bDNdlfCqKCcZdgObtP1weAKR6Tu7qMnjR7X3Q422oQE8N1SyqLoMXpfeG1t/T/5+k+7nXSD5A7blT4dLp2cte
Sc+l90xcSZCdSeIAxfBXHrDc87kTQZ7FyblToG6DvJpk0ZBpkcIJRICXNSBP8FkOVHGhR0zbKtLVJkmhOzYh6cnA7e97O6B9w/VXOdOCebSw3PO5E0Gexcm5U6Bug7ya
aP1zLtfFqWsTi8t+yQ6zesHkYeuXosApt7e7ou/pPi6zhX0cNWsF/WtZqxmWmos75XN1v39yRwxfzQH9c3mNwQE6VQgQXLh+sz+0T67Z8O3YaQZ83q5B6nYZLjYojIcW
CYxjDNCqge7yTMsyJV35LbDc87kTQZ7FyblToG6DvJqOcLWV4hlbobUpB9hG5opXb+wIxiTKXX0Ajc7eZIMkiuciDPTnZZazCr2nLu1ibwt5vWPfKQEpYfAfFkIoWwGD
xvrXe3MS6DVjYyQOUuooWo64hFGigmzSxv33v/XbSZUHNG/67ZZJi+WUBuZSWp+wBiBlp/lyq7Xh6LodLt7RPVUC1pF3NxVDS5rxnsHYE7i/lQs6W3xAGhV+3WI/bZhm
4zj43zB9ba19GOd5htp03GDpvb7r68q35y41tG5ECgBODxtqhJq/8EVizBD+xjqYW6QhxvmxAEEPBA5fMqI/+PmE0/THssovMK3o/4oSz9nFi5iCRQI1fX9c8gM7hiRG
1tLy8QikJaGPBj9wmyJ4bKw4HGns5yTPlrVLa51nHdw0kdaLOix2tEuYezhKONNt3BKQZp2EOrIWp6nImLFO8tqpJAfSvMlaYlKdHcks0XyG0j9W7wwlpjCqFvhZkCwU
g25GP2MC6c2a46jvnJbkf1Uh59ERS610z74PKFcPQiouccpQkrr8MiODFqt5gfrPQLfcNwWVyqlTPFJKx6pcOR2eG+U5t3hW1UPPlIpTghfnIgz052WWswq9py7tYm8L
vfsXqFavtQNAIEuAKJWJhEtoybDiruuML52iuyAaIJvnIgz052WWswq9py7tYm8LvfsXqFavtQNAIEuAKJWJhIRyvXa+Kzq2PDkUx3yY1bTaqSQH0rzJWmJSnR3JLNF8
YOm9vuvryrfnLjW0bkQKAEQbrHlWAFBTEcut+q1QJcTeyJCdg40YLR8y0th2HuBqjriEUaKCbNLG/fe/9dtJlf7jpIisLIAD8dNI5F/3MBd+j4z9NqSCJWA4a9STAAly
5yIM9OdllrMKvacu7WJvC737F6hWr7UDQCBLgCiViYRYFOCHs3CGuF7ZlZnusI33SW9NF6CKBuHLdrfZ8dEq9i+xKsp6fF0HcIXyWZhR7068KRIp8UkglqW4RoChjP9K
GbAc7AntPAxQ9pO4dUAJWvD1Ga78B8bdjzVYgNp1r9p0nbz8xlSO717b+L5SmK8uSW9NF6CKBuHLdrfZ8dEq9i+xKsp6fF0HcIXyWZhR707Sd/apBaBrxsxREpUIgQve
MV3DSXmD9zSEpIpSHEj8eX/hpoqEoKzZUrmj3ABtLTBUdXja64hp8q1sp/rjvLw7VSHn0RFLrXTPvg8oVw9CKlsLDZFr+pFseEz54gkbXyjYApdgYp9dLNyu85es2m3K
GbAc7AntPAxQ9pO4dUAJWvD1Ga78B8bdjzVYgNp1r9ogM22FHkucRPYeWu4bM0WAE095AXPrtUmkFmuFqMnPCo4R8zJhe3kc+ZAXe6nIBLZXLvl6RZcAL5GmgmKemzDp
JNhv61neDU9fOxEMY1rCqW0dJMul6zgeHMxKJ7hLkYohB6HIW05v4Gg5DJ8V2aApgEeb8SDsFbkp+aeRR/Q2uGx74GoJyO9XEjmz77yLuOGFKCornt9Rr3qpXzktqku8
GbAc7AntPAxQ9pO4dUAJWo4R8zJhe3kc+ZAXe6nIBLaT4RbMJ9ukgIDYJcZbW72ZnxQu/mKFxhO7k95f78sJr/D1Ga78B8bdjzVYgNp1r9ogM22FHkucRPYeWu4bM0WA
+RPug31UuHibMStN4gjZZ6w4HGns5yTPlrVLa51nHdzPEr6T8ipPD1hUVhDjcDZjlQILCgvjKdG97chbCSbt/WDGMh3/fb7gs3BPnj74joHKDtvmmCtlJ55g4xRBsiHA
MM06zAsD2tJ1Gn4dkASwNtKNr+ytxIWeCEvmewe0PrAn/C+g6xeNmLohy2/SLj4yyQURs9dieInI65AkphswgDxcQaQTE+KVzGnmsK/nudLaCJLycDlDBlH+WiQTW0d3
yijZh8LmwfiKibX/WkCyZEN8issZY3Du1lArmU+35HOxeB1aYBEhpzFZBeNRLDHJMV3DSXmD9zSEpIpSHEj8eVMUSXKO+kqBc/okKie1QKjk85MZ62NH1GpyZT9Rl6cN
af30p8u3P6Pp7E/RjvIh6DH/sh1M4vSO52NaabeekjYefL7hi3dV86z1sRh5dFiSqC8FN8TpnE/kVLIpmNKkJdzB8BKFr2BpXuw7M9aloNq8YaZI0Hh7OPDK7EI3VHEt
B3DSdK0byyrgr9R6ql23HKgvBTfE6ZxP5FSyKZjSpCWOGC1iuItrp+82pnO4DbX9EmQAIzEthck1lJ1KBnzrIWVQBlmLzNL2ISlCVY6pgPCUwSf/6d47+7B/DCLAGTKp
qC8FN8TpnE/kVLIpmNKkJcJ05p22ejztAxf2sCaErpx1MzF8cbppagb0EH15dCs8RRHPLWbYozHaqLUqktEbzsS57ye6W3pBOgZkPScYRRZM7qKKZA1oio73h1eKmdie
XysWvkUPPKsMjYcGvMYzNbiYfY7uzhqTe/2YwH/7RbU3qPw4brXWTNX4rxAYpmSQpw1jADsXK8XmDMHIZltOtgH/th2P7CBqU4ZBvpds7SVHPALF2ihMzR51Rr9pvweU
yyZ8LhZONv2XhWMO0lW+dp/ntXmEZs8SNiAVj7UC6+amaMvF4VMtJdYplmwaAySPVOtZWX881NCHQLyHUmoLg40AFa721l9nmOw8ZKVz95kDuAKPjzG0BxVDeJF8F/jb
wiL4acK9sN2h5/5Z7iEparKX/U7HTJCLIA9iG8RVXOl/soo4kQqoWMhM8vYUx9PRrt7cQRztH5QLVpqsf8lQLPgLIzdsrqZ6SrEuME5fU/l91DrU5LLqv0sVP4TwS899
8GNgkyrWLUMwvcMBAmoNZskR3Y+ub1UiyG7wf3xIlpkwkouibZ6F1NGdhddvP3VKyRHdj65vVSLIbvB/fEiWmdDkQ7QPOhXAg4Mfbglknpka44jErHH6VRg3+WakA7VE
3UbQpo8TLtU5P62C33kpDIsS5MGFVFM0VVjukxsFN4CdOCBp/NBwhz7MzyLOziVX5AHQTXIOmNd4kIzh7GKck68B5WivnmaikmOklYEMt1eyfOC05uZfv9ojk8c0gFf7
+NKwOVZDiQdb5kqAtjQAYo4LzwAFl/1TNGWdpRt0dRdbYMZgD8F87uk5CYeEH+1MYREUkbT0pc0v4Fp8HdCj0PIQpLncI76EffHDmw9XUIa3QeRbaph15s9gRSqOJljJ
dbx5ffwoUnGHgzyhOz5KLHiDPJEAxTr+MV9W/HzpdQnyl1leRLa46vuaK4KRppb861f3EbK0KIF0xNeK7LVkcGwE2aXjCKOtgGa9PbklZ4HDxrnCfeBPBQigbwt3Rwm1
WlkmP/lPdzdV6z2Yd0L7VGus1Pxw/gMncMh2IeVurDFzd2bMIk5y+b7hAFVDXxjaCzA1giAT9fiKUkIvtLOxqs7N3Kasiso3ENJF3Vq/2nbMeWPmcTwBMPWPo8mdXGwK
M80io7RcGOSERyLZKJy3r4fPnUocYhLdJQeboMcSy2lYFdHTkTzYmNhSzHmRU2hwnFrfxILA1+M1qJrrdRsONXN3ZswiTnL5vuEAVUNfGNoLMDWCIBP1+IpSQi+0s7Gq
+JASm+dUlAx/oyzeymRSdSSIgzcDwr2ws1adpqayikcxsUfkMkvKO8mmX6YN8HXiwJ3dvzgrmwJcq6wjFyxiqnRcGJALvthodQlGxlEtYdVon+bi3u6R+XwJMZ+t4Fxw
BStOHwZg8x9iM7M4icetBYW6pm/3vvUwCurvj/IIPkZpp9BfmRG0vLDcj3KXIr81dtOYatpnNIboiXichjmXl7Dc87kTQZ7FyblToG6DvJoSQjAK7gfnaakqetvTxYx+
yyEU+UfjHvM8uU/3G/OOWYgBRfQssOe7KAoIpr7/Bcqw3PO5E0Gexcm5U6Bug7yaSjijyNwRasvGnEAjcM0Wp5tGT29jxyF9lqWuJXJfMmhoOFj1zLCtLEw/kgSUqcbe
Lu3VpzBYA+WbRhplivSVFewG8dhyDv/KiN3U68iFvwIjzad4m9DbrP3Hpou5U6U/j3KOFvFLbCZ3MRPkQa7kGmM4OqppRoxgYC7VBkV6atx4l1hYxdWM8hglXgoWmacw
7HS6xhAP9NLizZ0i9nqE0I4LzwAFl/1TNGWdpRt0dRdbYMZgD8F87uk5CYeEH+1MDYBRsT4QUx6JgSWR+p7NiOTY3nIXmNyT7IqByiudxOu4W++uj2AvQyf9shkDROhV
zioiWg16mApuqj3kgOdwUhZ/WPs5g3QA5HcamPo/jKwl79J1ahE7cQjW5PXSRvNgFyOvvRHR2M1cEZ32SbW+Etvv7scPSTMdjiRWUzSHI3Mmmm3ITT5Sri6eVw107DdN
MhaXjZtqbNWNAySaFuzaDmLtYTQzTHJtCLesKuUquMyw27DseU4sD37CTI6D63v5Ng/+ENDwpy0XQyP1JegYT7+PXGzNFhoPXGsrpJtNdccxnye/fhk2Rq8gZsXFvBbk
Ax+ty6+KVLbt1A4gGgChDrWRhuChANdQ9KdTcSZytlXCMaszjrWuylRdfmN3xYrFU87LEw5ouHjxmBJ8FDHTbvmpYRmZf1HuGfO5MrWgHUybs5SnKqv2qN9897bs7HoC
zZeyNVFOovor4HV7Z81zYXmvSsEIhEVhawjMUP2cjlQkBXsg29haCoHUlbmK/n0gnRu+6k9KS/9uQT10PQ6gcooXWrSN+MhWs18kdnblMlnjIezt+EFYhHa5b/smJ99D
zTjF7Hq1vjXUFkGhieoktGXdtqc/ef3hJI0MlpXB6CkqMWnGd3Sw3nwYvBKcf4xsTCH2dhdy3Zj7I36Sk0/YRmJu4OJ43r/pgsYnaHd3zJIWaR+4BfKIBH39aLUmg3SM
Lctn5/jrN/l2tVLGOKm+9WjIIpFvWYVZacbpx8vx8ceZfCP/XvWbfT5dcLY1dh1Wyzzw7W+o+6l0ocHXkxl9DXO+011YpGK1x6hsFc2dMVgBxO8XyDCigwqYoCu/mbTw
gtZan+Zv0dRzL52loOgT1CQ9al3EBjnOGmR74zIOPCJj0NzDYsp2RLdi94WIpWKRHlBzl586tzQeUagl27WfRlo/HJmnVyUz4SKyN4cmfztsSlZVR+Hg1tQIdUf7wmDu
qsfloDQpsHdUF8xaeWTPPIyjPlFf/yeOQIPCnGirsG05dQw9FwihahZwsbD0ZsJfpC2WC+rken9jA5fw0Tn6eY5/KiK0dM7bf7ergetnat45RBM4yPmZ+AmlPsxLjlOo
8JoSnAHWaUwuSVzn5GP6JLBjYIA5M8EHcSPlSvuqEpBxQVnaDR5XaZ4sfQI3j500ZJCoIfK78yP8enlVTxD0j7Pqzge+g22Bp+dJaQJvBsAKx5nfTZ9ni8au/H5bvlVH
u1xdSfuiAjlxdkyJtp52se4FFNZ/2Gb2RS8RCvS1WuFG96iCYn/rexjm+Ou4HpWwhBPOXSK1ArtQVcC6yo/Ss/UPz/PbpDbwwEJeeJaxDev3rUqOOiTSIdhTIMg5HViu
YrQbBGEIsMZyirwI42iOCHsUJQ70k7Me0Mq/eJmyjzI1+6ngS1UPmjnQODUwjp7+U6Me7iisvZ3IezuJClkkw8x6Xa3g4XmKGi/ko9evN2LSnEc+Pba0aKAAHIFrJR8K
Uu7B73QIikzIEvN1L9W/qNwo8FNwLgmRcBOo7MPJKgKsvmMHxZ++1x4DCg0pRMaNSyIu35ryxKO0m7jdzKb0LlPOyxMOaLh48ZgSfBQx025abiWGvqawvVvtqOGi/n69
m7OUpyqr9qjffPe27Ox6As2XsjVRTqL6K+B1e2fNc2F5r0rBCIRFYWsIzFD9nI5UI9NZiAwrge+VLCcWQJ+d2p0bvupPSkv/bkE9dD0OoHKKF1q0jfjIVrNfJHZ25TJZ
ITLbSOS6fIIzUBjJ+ZzjKc04xex6tb411BZBoYnqJLRl3banP3n94SSNDJaVwegpKjFpxnd0sN58GLwSnH+MbCciEaVWYIRS16b1ob3yQMxibuDieN6/6YLGJ2h3d8yS
FmkfuAXyiAR9/Wi1JoN0jPnmerGR0MHXHDRQeP8rNployCKRb1mFWWnG6cfL8fHHmXwj/171m30+XXC2NXYdVqnOLTD3GE5nY4rhSZqVGvdzvtNdWKRitceobBXNnTFY
AcTvF8gwooMKmKArv5m08ILWWp/mb9HUcy+dpaDoE9RvsgNL++bkD1atIH2p0PwMY9Dcw2LKdkS3YveFiKVikR5Qc5efOrc0HlGoJdu1n0Z29699e4N/9KJ+HLRZkriy
bEpWVUfh4NbUCHVH+8Jg7qrH5aA0KbB3VBfMWnlkzzyMoz5RX/8njkCDwpxoq7BtZC9IGfWrVF0wfSNlT3cBHqQtlgvq5Hp/YwOX8NE5+nmOfyoitHTO23+3q4HrZ2re
af7DggQcmaiYK7AfT5hvofCaEpwB1mlMLklc5+Rj+iSwY2CAOTPBB3Ej5Ur7qhKQLXFZptCUdj4NUXQPRtYlMywL27Ry6VlTMtOTvHBAn9+z6s4HvoNtgafnSWkCbwbA
TPlXRgp9PJnHxKjQCbgPEI7yYGgNvtxGubaZJZH7w+Nc87IOTcgLSaToZt+lYHjUUHIZk/aT4ArOiIJSUGSJmLbsLVe06vnrUpRWU0DJUa+uyCcH3NKNi54OjWYgXTg5
uUan0bLJVdQiXf1g0iTA47aoHQeU9zZ7+RvFXBPWg4LLSUMflfB58j/wHLad7VLbCY1Jz6GikyAl7rhG2W/Q4B5Qc5efOrc0HlGoJdu1n0YGkwa8VIX7iJjj2pui5jiC
bEpWVUfh4NbUCHVH+8Jg7lO0kwjuKmtr0vTbSm80KyDAcUATREv1NDlmylocI2QH4BXXffItfpenlpC7GzKbaLM/EN+6bFB2Rj/+sDF4FyrzLJup3x/2Z+xjdyymrXEE
3EVrZG5BNiHdyJhAe6k6rbirAHWZbueqmGEC7TtuYOc1cAtgBy8tF7C5Q2jX8y13Xs1XrYP+se5JkWQNtxqAg+nOGQxDHQ5RoFsxZr59YiR1hzdDo8JIkIYxe5iFpulp
a/vOvf7PFwe6d2Doi7e2cbPqzge+g22Bp+dJaQJvBsAKx5nfTZ9ni8au/H5bvlVH1wHE1jkwrb2y5cL0y/9KzO4FFNZ/2Gb2RS8RCvS1WuFG96iCYn/rexjm+Ou4HpWw
cUFZ2g0eV2meLH0CN4+dNPUPz/PbpDbwwEJeeJaxDev3rUqOOiTSIdhTIMg5HViuYrQbBGEIsMZyirwI42iOCBAUAwm9xW6vvEumUWnB+RI1+6ngS1UPmjnQODUwjp7+
U6Me7iisvZ3IezuJClkkw0/sLPrIMwNJHspFMK8TXebSnEc+Pba0aKAAHIFrJR8KUu7B73QIikzIEvN1L9W/qNwo8FNwLgmRcBOo7MPJKgLdSlNNk+ni9y/QrsYAp6V+
SyIu35ryxKO0m7jdzKb0LlPOyxMOaLh48ZgSfBQx024Ci19b1qcHqLsDgUswehCam7OUpyqr9qjffPe27Ox6As2XsjVRTqL6K+B1e2fNc2F5r0rBCIRFYWsIzFD9nI5U
ePTEdmsbKcXX2wcVp9hJ2J0bvupPSkv/bkE9dD0OoHKKF1q0jfjIVrNfJHZ25TJZjrhUyhV7mJp6uTihYvpQdM04xex6tb411BZBoYnqJLRl3banP3n94SSNDJaVwegp
pNQc8e0MURdNomo0+98oGUwh9nYXct2Y+yN+kpNP2EZibuDieN6/6YLGJ2h3d8ySFmkfuAXyiAR9/Wi1JoN0jBTIckXs0NtcjBNCNGDLf/xoyCKRb1mFWWnG6cfL8fHH
mXwj/171m30+XXC2NXYdVs1nfbbiUnVwa9jrHROD92pzvtNdWKRitceobBXNnTFYAcTvF8gwooMKmKArv5m08ILWWp/mb9HUcy+dpaDoE9S8BEz80USo4bS2s8M72+MB
Y9Dcw2LKdkS3YveFiKVikR5Qc5efOrc0HlGoJdu1n0YefKbOZLRVu7Zx9DMpZQ5mbEpWVUfh4NbUCHVH+8Jg7qrH5aA0KbB3VBfMWnlkzzyMoz5RX/8njkCDwpxoq7Bt
tfe7fMlnp5T5STPlRF+c0aQtlgvq5Hp/YwOX8NE5+nmOfyoitHTO23+3q4HrZ2reu/cZaXD+ylCv7EvQOxs/ZvCaEpwB1mlMLklc5+Rj+iSwY2CAOTPBB3Ej5Ur7qhKQ
cUFZ2g0eV2meLH0CN4+dNG/TXcuaxpCl+hx3cMDWrUWz6s4HvoNtgafnSWkCbwbACseZ302fZ4vGrvx+W75VR9VdCNRQyAoy2TNcFNS4/9juBRTWf9hm9kUvEQr0tVrh
RveogmJ/63sY5vjruB6VsHWHN0OjwkiQhjF7mIWm6WlRUGwO5lczag5UmaAL+wK4961Kjjok0iHYUyDIOR1YrmK0GwRhCLDGcoq8CONojggaE3BzrzZrqgZysx0C4u/v
Nfup4EtVD5o50Dg1MI6e/lOjHu4orL2dyHs7iQpZJMNERvAhIDLdYQXLL5mwNDCn0pxHPj22tGigAByBayUfClLuwe90CIpMyBLzdS/Vv6jcKPBTcC4JkXATqOzDySoC
h7cj3dFfja3lSrVbnwr7hEsiLt+a8sSjtJu43cym9C5TzssTDmi4ePGYEnwUMdNuHlYctV/2YDu76jL2FLoDzZuzlKcqq/ao33z3tuzsegLNl7I1UU6i+ivgdXtnzXNh
ea9KwQiERWFrCMxQ/ZyOVIwe4/3myeD/UKJfOwT1t8ydG77qT0pL/25BPXQ9DqByihdatI34yFazXyR2duUyWc4/f4ZsYICeHOYHqtrrgCXNOMXserW+NdQWQaGJ6iS0
Zd22pz95/eEkjQyWlcHoKaTUHPHtDFEXTaJqNPvfKBmAKz522lnNE2ZYezBOCqfZYm7g4njev+mCxidod3fMkpvsE8kP0I8jm5ONQqJgAuxGJiienFNKIt+UXUiZ3XST
aMgikW9ZhVlpxunHy/Hxx6+DQUjXHjJKHdGSAJAd0FVxQVnaDR5XaZ4sfQI3j500uiqhS3pL+5zF4BwJqHYYTSBw9xtSzHU7yOxb2K1a2PyexiR9aNiMr1BAP6qOy3LN
2/bKtlshAIdjfLyduhFtRmkH/K/6HsXNNKyc3iQknIPouJnmKs4NK40F3qv8wykTN+iBRBLEwRzu8/IGCiTL56ZQmUtpZDgvVDkLncgar0/+N28FQ4YIqPI07RanjE1A
D3IJ06nQlnYSsVPNWvD2YZl8I/9e9Zt9Pl1wtjV2HVYomCj1WzxM4eXXrwmLCYC2c77TXVikYrXHqGwVzZ0xWAHE7xfIMKKDCpigK7+ZtPBtIexqvVKue3w34uMG8ZGR
nRu+6k9KS/9uQT10PQ6gcpuWjHvWbCoz7rFlhsyPiS/sdzOOynP/M53pSLmT5qEPg7nIJjEnQimcYOmRF65dX25p/fmGqi5f9yuET/1k5Kk3DlfZ2XtWSw1Rit3m8K30
2qkkB9K8yVpiUp0dySzRfG5p/fmGqi5f9yuET/1k5KlspHrLrn7OZd645CrxwvmIsGcMTDxpvINECDkaC9Bx+etp2Po0oUFNVy6BPT0rJ2LEQ5WRLAZ6l5D/My54STly
Lbqrj/1tduI0JTBC+RqS8OcgQpYRuD5YllP7eHdrRhUM0Kr/uZmSMIjahN8ZHLMuKoktvUhZCOdXWnrvFScks0sN+BgbbglMoGBi/oPY5oWSV4VENM40f2sSeXIg+W6g
+YmR8AE05iJWeeJd4Zpm+673Is5OTCMqNWYuhjHjVbn4/K+0oHq/POiTVP6Aa9MDxB+N9kJbIgOq2e7QJ7OUwr0jRkL178pl7vrxsFLhRcAox8NzTJKSAfJhkz/I+txP
iaOcvcN/oWkPf0n+pRp/Vy1ZJnYR83s15d4MFW6GocncUkntkpYiJgS30ItvGgbYDFB+7PF58QCULK/1vCgZW3KNwfPwGwmen/+Lpcvilgj57s8r5xEUKs/3wJm8A1Q0
kfjDwruOxplRcgtJx0gnLfjWS+5KwMYLtqsu7CE2/oeEo3RJbrLrRlK2TltPtngXDW3iry758mTmz8eX70BaiNJL0f+eUGt8rD3jMkgvzA9QYytiHG2PlkYDpfh9kURw
CihTo9x8dc2nzHlsQot1YgnjtF1PbbSL3ABepSJy9VqCr4p4DfOxAVUmyx+46IswmGNGe8pl6mUZpSlgK24/Fs32YmyQMAWP2Z2LF7Qg/NGyBc1IJbtfov/rqIbxLKH7
nOJ2q8c2KqnO5pGQiHeDGgFMSW+Av9iwqsB9Ou/9tm0MUH7s8XnxAJQsr/W8KBlbC2rIi40uw4GLUXKjsoUdLlW1RSytyEkPvyW9FRZctC5wo0vbEfHiGDdvpb98wp/J
h4JZ983eNhpMApHfa787Q/eEPBi7xIGv2zgV6cX7CESnrnQ67YLWQiWFzXCRPbbWPKDbHxJHHbfeRzIr5W1Ys4doqEbd8gx/YKvVnG8alKrUefHv0bdNUVt0jjzlAetH
Yl8EqqTTnx+JY/A7hsZkEKqaDIEn01S4utfqdfhWOLyzTd54Ywk/CnnhnNQ7a9a4Yl8EqqTTnx+JY/A7hsZkEJnypBtA68zbqAZZdyaZ9ttlFD6ro+ea82qzBX8UPpxJ
g7nIJjEnQimcYOmRF65dX4V3WapRMZ7CVulcsAo1RWvksLizAupqzo6ufK8Lbmgv15bU/A8ziT/TwS++vFSVFgkZxC3BbjUT4qYtzt+ooH90JG7zoTE4DchGvzKx73/L
6n7Xx7fb2sjJe1RJe9ud1wwokXyLKmuwoSV37jr2myCZgn6Ot/jI36ZhfLDhVh2aoZGyir4JyqaOZN6+BTfgP7dusDuac25EReEQDWYhyKW2OOVNBrGwEZTIsiLMFOw5
VC3dHlx9A9mxoxwDyqFujfOg8s/aHY9huDXV0u3r/ykN9X72ZE48j/ftvXPKV6x0ZTeNJ3EltKHrY06VZ2g4zsIi+GnCvbDdoef+We4hKWowp1vVpF4y0bCJesqxD/ds
R+XQ17yVciFn0teu1gfDn/iotzioKtZNxYy8MX9CHQ18KABJgcEUIo3cT/pNI1cKYuL3AY9GBvvibSh7aIvghV/6zLDfoPfkVKfnOhaH5X86tfV+XH9E5WtRTgyu/3dF
9SBEX7jeFqhzYVGT58gP4xBBQdcJuys5/FK2gEEcfjeVwsb+uPR2lyApV1QwTYlIyOtUElWTz5N7xL3TP4yTyxrjiMSscfpVGDf5ZqQDtUTMvSbL2iGAwErsqGNac26h
NDS8sYJ+gPq9vFfJWlQ3SsVd5IaYNaS3aJbAX9ZIY2OrAXMLBlCNpfgmF/Bj4hbNB0iux8rUoJvPwElRkubF9ibHbg7Akm1H4E8T3IFl97XeXekzfgGvJ3jLDQv/XvAb
hznndkNp1wU9/YiOZJ8urCAHxV4w42/CGkuvd/kkXcZ/0Y1I7kiR33CUGXUwz7asv7DQt6ie4pqWc8Tiuq+RRrxTqOWQwIUD8K5b3Zc5jQ7Wn1rCVqUx6Lvo55zqomyV
Id1FdkF9Y2f26tjA3RH1vB7SS2uCwgZP0KSay+QnUSHbeV8OerGFziCtFyhB2BwMz97IqqdV6WekZRgynbXqOrtAOxFdW3Y9EqFfSMpoyAgQIhAFvl6Ui/6dE3IvwPXK
8cs7oLqheoeYmmTyPZ/T6Pk0s5LfYXTxpuXgzWQEhkwFK04fBmDzH2IzsziJx60Fys5+d1LWLIUzk8A4UjJClFftSvq7FRlzoaCDJGC5r6ZJHqg2Na+sri+0S+ndkqpN
GAZesYqrkxou9YGmspGhH0/0HaNDInWP9uAPlxkq4kPVcbHybk+59QlQzlMkuGb7+loLn5Dpjrl+dTqsEgEcmNVxsfJuT7n1CVDOUyS4ZvtwWjwCBY4H6cnovPLVCXqu
u0A7EV1bdj0SoV9IymjICGrhBI4BQT78tp/ZrNMmIJ4CkImqeM1C2hN3uzTxjhC5RXe0Eb28H6nl3twsbxjWxLtAOxFdW3Y9EqFfSMpoyAhqbqUhPexmecusz7OKjM42
72qocTOJgMC7M2GlFqcVE09YKziAbWW1a7gmqZ9YK9d+26S7lX/7K7RwzMJ3rg8+CJwL3yI2oXIWE/vNov5BtxYYx6sv3IoDys9cnLS1JjuU2VIwjw6TFq9V11Zxkcu2
gB2OQzVk0Mc5OLbZA75WeHdb534wsRvANH/asxzJrHxYYF2p6pko29LBgeNR9t8KuzC29FwvVlIqyy+etodH/M9ry6rg7+lv7ZcsdG6SYL2n3gizQPcPOdcTS+gTOmKJ
4+kAT1Mo5kl7lJTywyKvEeFLm5ztLvzL/b99qlUz+rv7DxEs/66L2bfmU6RVY6nG8ShLsRHMnsdhFqBPzzjaZXEHFErppmd2Lz2lv+fbEYiR4gFIKJP1BryF2iFu7loS
rzAgRISBJqM/LN8EZgI5nVefqf+sbIkmVxfGkZ3x/F+nVtu5fkaV2/Sn7sna6ZRoVSqQGZlc/bvFQ+llt7ksgd8OilRorXociBySVt6t4N3dVN5PqzvXteXuPVTCnCPg
rphHOrHbXy/Kk3SSJXDd9WbLX+YGeR/et1wQ0YjvkjuccYNJqPWEBUaXrkLPYgDUBeF8XNzfnwA/e+Pub/An2JFe/YwPqdQFSCZvxIS0wC9AWBUAT8N0LBOmQ5OsLdu5
kFcwl2bjuxsGVfN/BVcS0Dx3RRmHV+USIk9rFVecRwnZ7Po0klzcD/dAYZKPLkIEjXpN72IJak3HOdBUjakfReFLm5ztLvzL/b99qlUz+rtIdGeihMaSIjNEKYtZjAp0
gB2OQzVk0Mc5OLbZA75WeBXgVKWO6du9E/YUjqb+ZdbRTUGesw80dTl+xX6dIqUe2Vir1qCck0ZEEkXieQ1Sza8wIESEgSajPyzfBGYCOZ2XUbhIwPW24eJJx7RyV5Xm
KJrenAdUn5TMFkz8lz3Hw7LhoGOLpatml9mCgyzNYSPTIsB9tOhYjl4VwOSWVidUM8yJTmVaqPZCgJnKNeai6HHglfIwTHiE+btfmrJFrIk//L+PwzHOIYxMhT/u+2mf
gB2OQzVk0Mc5OLbZA75WeAVVqs3nGGqoCkCzyasFXrEaKp1lffdU5XAHnHQ+Uw+6OphwATLtaA5C0EoIoK1V9P98zOyLVIGGcRq6Mr+q7p0BNLdP4Kh/mIcrMndGdL7E
w04ZNB0m27sv0riZEJG8aR7z1MqgK2vuwF4Cbzn8P7LIVeqrava89a5RAPzd96SfWtXKLUf+4eSugyEmx521hdlYq9agnJNGRBJF4nkNUs36xyX6F2VvFprt1yjkgPnz
+ciZxQC5pMsZPbMG4ecguQ5BKiefJkktYqlS6mDM17qopDvF0PAW+/Jc3ng52UPL7uX3MeDohZ/UzWUxu6/2TgE0t0/gqH+Yhysyd0Z0vsTDThk0HSbbuy/SuJkQkbxp
Ekxu0jQeY6k+RqAFSR4bAMhV6qtq9rz1rlEA/N33pJ8aEqmnEIkO4cBotuVx6LAM2Vir1qCck0ZEEkXieQ1SzfrHJfoXZW8Wmu3XKOSA+fNm33ydg1J9QdPmCSsoj4ky
U6bgO2hzpVM70iDAxRsbWz2UHhRP5OuAUuUz9JhC5sBWOj+QDZEQ6xunjVraFWF7fdj+SB6QfBXVBoQukfy6wiYrHYHHYPcbMqxytDl9gXLWjw+XAyK0VB0/bjMAmj0/
NIsDYZMCOUXCtdRl+rfui9LChFE27jFfHxHSGOWT+ldJb00XoIoG4ct2t9nx0Sr2dRfQzQe7PWf/YVqFuC2s5/I16SvxQEDX3q8i0a1Un6PISVW+ffuvOyJqDhT4FCAO
dm8aR3400lRy0X9yOnEsaBxeR/J5goMFZjwdPIsjsUFoaDSd+r09xZ/6JYfs7Kpjasae0SrPPqIUlNfLNFxMwPkX3myxdzPMfW/bX2ncBg41MdPRizeYTjWeYDeVmlnL
FPXoKFU5gdLT6RE8f5xpj2tkD+vshh0vTs19n8gj1L31n2yI9jzkUQq4AxtbQxbebAfQr7LGlyrljTRXkyRK+uf+SYpnnR5NzCAmOpPT+/9e2AlvuVNM1qHA9H/nAuXN
Tmiq2iUimcCJfv3Ek4A7tu+YE9V4904xDG34ICmaflIrFM6Xob7XPZDlvZHkOHdc4rff6aK2gF1OqpTbmaxyyMfLaKByphJ0nJebyikoKd5YPAcrhfVqRx2PB5gdGe0X
a7eABL4lxZqMJHlxyZA7W0WnSOmgEJHtFMuldaEK5/2PYm289KnPSk7GhmfTGUAVXtgJb7lTTNahwPR/5wLlzU5oqtolIpnAiX79xJOAO7ZVkFNnYmWnD/3I9qBc/LJR
j0M1LZfCtamifyNpbza+eZ77t4Lss+XV9IfJeoxFtfIrFM6Xob7XPZDlvZHkOHdc4rff6aK2gF1OqpTbmaxyyO/uQW5DPQYEc0o6PzBKqtnISVW+ffuvOyJqDhT4FCAO
dm8aR3400lRy0X9yOnEsaDo+DMKncFDdAJCE8e65Yz2u7UEgvYHH00gs4ev+/0ILnbs0VUmU5RSFkO9U0YfUvITlv+6lqZRDuGon3/uGUFZ1Iy2ysaKS8d5K3pNuN41t
KxTOl6G+1z2Q5b2R5Dh3XOK33+mitoBdTqqU25mscsjV0u89wPk4w+x9udheGxe4z1NJ/9+3zY2UjGFMVuZC2y6EhHioCVpyDJbCWzyHC2XISVW+ffuvOyJqDhT4FCAO
dm8aR3400lRy0X9yOnEsaMZcQlPtp2G6m6m+wo652X+RJARM/Hk+I4NzMAFUmx5HRadI6aAQke0Uy6V1oQrn/f2ExJK9ZPW2w7LkoydYggnNhSLDBm1bdjVpGwwWkk7Q
TkvbjECqyHfxR71N0VGfR4vTfrTLSqst0XcFv2JHOd5DAU+IhlzUKiEwGOfeSbWGyElVvn37rzsiag4U+BQgDnZvGkd+NNJUctF/cjpxLGgPaapyYQr05clfms9lkQKm
kjkHnDPbr9tNzgRHJGjlFCIW3rEfziDcxImu+sI9hB6VPJErA6zJaxSd9xM9fSf6T79jZcbf97PBlsoX4ec8sfCdiUmaYxfkM8UifXUxmcBnGSTpH92WT02mswLueNso
RK6q0VoLiyzL4hM5mmYYx5J3IcdZJJP7ahnMBLGbSRkkjYbJ3lq45+qHC55nk2Kf2qkkB9K8yVpiUp0dySzRfFZ1XgBzxhoOecFJFfYVDR4cbtwSHn2WUTxv4d7Atm65
cJ+aq+sCAM6H/ymsq6YsDQicC98iNqFyFhP7zaL+Qbc3PxnIhG4enjXApC/sLJzbWtXKLUf+4eSugyEmx521hdqpJAfSvMlaYlKdHcks0XxWdV4Ac8YaDnnBSRX2FQ0e
HG7cEh59llE8b+HewLZuuYKYLjIlnaLUJwby00mISghWdV4Ac8YaDnnBSRX2FQ0eHG7cEh59llE8b+HewLZuuX7CqLDfs4SknKaO6KboyxAj/JAIwXXYtrjfQ2TlDxpx
KUQ4MOY8TOL4inlOOB2rQzTla9R7a1gzpBbiSTQo7OqfFC7+YoXGE7uT3l/vywmv1o8PlwMitFQdP24zAJo9PzSLA2GTAjlFwrXUZfq37ou2iJX5+xcDObbxFJWgAatA
I/yQCMF12La430Nk5Q8acSlEODDmPEzi+Ip5Tjgdq0M05WvUe2tYM6QW4kk0KOzqzxTBF1x9fYS+VorD4B9MjdaPD5cDIrRUHT9uMwCaPT80iwNhkwI5RcK11GX6t+6L
0+ORcIRuMLiA0STwwoYKtC+FP7VOozjwOK+PO0NHsJGDucgmMSdCKZxg6ZEXrl1fVnVeAHPGGg55wUkV9hUNHhxu3BIefZZRPG/h3sC2brnRFQhlTHhzH9IFz5bdkr9C
DIRsLidBGNrOXJwMl2QYd6JImbzO9LDNZGsv/EMA/LvPvI7vhHrGIr4z8fZCz1Uh4+taetYylgUMRkTxOm2tOrMxvIL9R8kq71OuGA5B1Gfk6kqwZqUrYUzTCsvraI0G
zSU+SAcAXhiVU6sk91xVrqJImbzO9LDNZGsv/EMA/LvFhBTTE/zLgtgfxKcUIqrdJ8OUB2v7AbjvlwZk1T/PFE3kprhZn/RGw+XSlpGPRVcInAvfIjahchYT+82i/kG3
Nz8ZyIRuHp41wKQv7Cyc2zVPy/Q1RBAoATpzeBOjcc3iKR/gnObezTg8WbSr1Med74727CC1fLkIYMJuxBC73a4s76+Tkz0WkmsSkzlyr/EMGFCcZk+MX1dyGUiO8/wJ
+RPug31UuHibMStN4gjZZ+Zc1P4NCo/ykdIfD8cAjKpErqrRWguLLMviEzmaZhjHknchx1kkk/tqGcwEsZtJGYTmHWerBlt9zxDNkOHg4z4xXcNJeYP3NISkilIcSPx5
eDy8fzrBEWgWnXeBxcAxtb9MexTOziCEouZ+kkC59YuVwsb+uPR2lyApV1QwTYlISkkdhaRRDe/v+MkFeHUquysd96uzpCKGJUGJWHnAzpSWlf2N6lXDvwVmgCsPGLCT
VOtZWX881NCHQLyHUmoLg5Zhtdc3C49K/Vut0dQurnGGd3vpSumiCB5abZKeZgabKgYr3uoFME/O8vsR15qSIi26q4/9bXbiNCUwQvkakvASZOBcBsV4S3Zvg5Vjnd1O
KChz+FrgxKVYzZ+uTjULNfIlvm/HKjqYUMTWAm+mtJPUJy66FSKqpKkQn5j2fqnSavSVBA7DV1FHwRHrx5PUR3mcbQOrZFWvCiI/pWNRlsxmAwMwaaYCUlptZ+PduyKa
p650Ou2C1kIlhc1wkT221vyBJmIcvBRKa8UY7Vp3shxJSnqlMQQlwxyAk/Kb6Z9U2qkkB9K8yVpiUp0dySzRfIV3WapRMZ7CVulcsAo1RWt6woSDibZlb/ZgYfk3b6NY
O5pvdnVdg0cUcJFO2POIRlcj5jPNV3LFNuhsfvcUHAV4PLx/OsERaBadd4HFwDG1tpgnM3ZSMLTvNIzSpRxxsIOR7WliRHpLVBiKQSgdWJKCNrg9JL0e5Z1rQ9W98LkV
4V7S3kUcmsYwkEfd/j4+Ycvz6Tsi1phekOA8HNk2b82PMBf+ibriWXwthZR5IH8cLQ0e3V2qtyIKB4VS02oGreQB0E1yDpjXeJCM4exinJNKSR2FpFEN7+/4yQV4dSq7
Kx33q7OkIoYlQYlYecDOlMBbb9kM+8KlSx1lkX6HekqBJjdHjh2gpm4NA1i7RS4iGU8wjUaCTK3VQn/2ikp01AhH7srfaybXVAhw5ldLOhp4PLx/OsERaBadd4HFwDG1
nEGEHnfj3veOl+6z77BHD25ZlgSl8dtqnYWyLt5rcKvuQOikC+pPEptA4bP8tlqgM3kbhGlBOZUyeLky0ZPuXM4qIloNepgKbqo95IDncFI43c9Yj2ayzyk7r7tfmGCd
nsX/9aR1g0A7m7eQFfHUhDBZ78nuxuQfQT47mzmvaxlrwgnf5Ga6rBGU50POnQN4zso2l+ltyoZ+fDp+FMPrJ2+D0MzaH2dSOIl2Q1P5Z6yAQYEru2pnCwOp6npMI0MX
lJdfru7le2EPwAlAvj8HCxIxgKnVbCw0NbEMgJLCtslpAkERB8COioWzYqLkP7cZCzjWlOPtEuGsP6wjDRQhq2DF1aqd9flzc9rabd0BwfwbX+469DnS50B8CPdwzLqi
zQqAtGVpHiuR89uS/0GcSucrnusb83fv5TEl0cmw/BoA1nlTEmqMu8hNJUDGZ5Vm0yLAfbToWI5eFcDkllYnVB9irc+PCXxtAhIB3jdEN3SKQx20UiX0lq4mBesM9yg9
el1mzA+qlbXOvjlBPac74xGQ3BHghU53p5aPhgTP4FgxikWQ0JFi0u9kRTfjtBLblIvQtGn38ctrT9Dk2a01a3T4OJhK6ee1gyH0f6NGAEjlPG6Jgii6rtSFVT0VH2oV
8iW+b8cqOphQxNYCb6a0k/v3LniFuwqa9aa5jOd+gPB0JG7zoTE4DchGvzKx73/LN7PCaLI4cRjhIL3vgwtecpSL0LRp9/HLa0/Q5NmtNWts+BBrwJHv5MvO9wem9BXk
5TxuiYIouq7UhVU9FR9qFd57J561U4oT2RM+n0mBkunzb8do/66j4UrTDXlOnxibIpbgsLsscCcy6o3KaQ692539l5NS/3v383W2sq/yuXsxXcNJeYP3NISkilIcSPx5
rAC36jz6WE0HG+/6C0E65LkcuMTDlrRWqEhVSYKTRN+3brA7mnNuREXhEA1mIcil/bFon+L032VyjZi5FWJglJXCxv649HaXIClXVDBNiUhioFpFxS4PIcl1oKs6M1bn
MjhY8LsEnVchnXTyBSFIVOqJHmiBrQ0wFwvhiTtOF3CQ8Lj2OgzrTJX3UXR6r4Ak5AHQTXIOmNd4kIzh7GKckzSpd54AIkMsKkQX2OdIql1bpCHG+bEAQQ8EDl8yoj/4
pMyqgotl9U8jhvjpyarO5/pejV6aZGihgyJki9SqrOM2/KHVzILmIEDeE/XqWaY6jgvPAAWX/VM0ZZ2lG3R1F/WcNVHBBBg88s4kZ/meGa/0oDwF1j+xPHnXQs/BPM56
Eu9QA/zwm/lcukabo7u5Y3ZU4RymqzXKguwaUlBgoAcPgFbNOmGRnkwnJBDiQ0vZ/sKl2RZR73owYcmaNAQfHSLTPin9jplCiVD+XBlD90dVM/J9o59YjrbJgD48Vn2U
qnX7OUNP+4IjZjXkF57DSlTGSAvwej4M8UJF1QY7JEoGZK2hnmAdyUViB4tPv3uQLoSEeKgJWnIMlsJbPIcLZaQtlgvq5Hp/YwOX8NE5+nmOfyoitHTO23+3q4HrZ2re
FuIccOgx2LZs6m7rEnz+wIDt30qfGoYxDvQ+fp0vTz3JeWaEgIR2KzYM6+p+4txnXTRj139g7yvxfVMItO8P3goLlPJa8RgRKalOD7Ro8QbASMnND6+C6gntogF8RIYC
3rs0Lzkong5HsRvc28VyTrBjYIA5M8EHcSPlSvuqEpBxQVnaDR5XaZ4sfQI3j500I1IAhhTWmjqzs42Qst93PxTgAH8ymZeKYQGZCQPAtCN+D+EoCm5UQwjU0ir52AQr
fSI4GUiSDg/cT3vbODBDK/Hxqz/31rHlw+t0TT+cp54PY8sSqUwff3URBC0NwKRCHELCW2M42m+VgHAiV31Hjh5Qc5efOrc0HlGoJdu1n0bxppkcc3qI+wXYeFs5oXj0
jthdrsVDm9KyXQ2lF1LlN28bE1Lr5zrHEcQ4w+qqGW8URigqznjYzNTCW/lJwlTYhVWZCPBt9cp79A5V5P01wnIN2IQQqrAc1/jR7WkyUp7i0RGSroq/E/WlqBNchxjQ
qsfloDQpsHdUF8xaeWTPPIyjPlFf/yeOQIPCnGirsG3KxVVdQS6V6nebgVeM2y4Us3KrD9rEXYgyRjLXghAujCDGWLxSlduWHwiWXsWr0gOON9goCQNlL5tHu/37Ttk+
9964RQg6QKRpYsQvlK9mXEhQ43V/Eziz61QBeKEwk3iErygOa3o7So+NpkxldU2UmXwj/171m30+XXC2NXYdVss88O1vqPupdKHB15MZfQ0KotMSor7jioF9GrMY8fxs
SADFI6Ez5wBLo0FQ+NEGJVJPXKHT2d1+8piBMgyr5YlhVnRWKf5UgOwkh6JVLPSYuz5PpwNw1InNx6nMixoYXqUYZCGoRFkkmK1LubOuAuoBxO8XyDCigwqYoCu/mbTw
gtZan+Zv0dRzL52loOgT1CQ9al3EBjnOGmR74zIOPCLrVNZsDxzwcGJP9O+tEJ7wYlH3zz/0aRaWCKSMbV9xLAthPorn7/DLBN2+8xCZViBnKdf1xrnCYrdqkBUeDgN6
wPpNGcSQtUTWBhaPWycar+iBe47Q8EHSCYNRxRmuVi1l3banP3n94SSNDJaVwegppNQc8e0MURdNomo0+98oGZQ+cGrNxAzy08h1c5mmyCrceU4z0jCMTzAjMdzqsAaR
k5fM+i5eU4qQqwYz7v4kRnJGlgEQNJlSZevWl5GWjUVKP/IRBkPm7/MH4LxzpbIDyf1PjaDqbW+C/C/gDh8krWJu4OJ43r/pgsYnaHd3zJIWaR+4BfKIBH39aLUmg3SM
GailE6k2pnINkf9E636Hn2NmgWhxdLsyzpQEzo8Yi3x7UVC9pXpWXOeZmSwCOldJpypmoox6q4B8zGtH+n9XNXMNxBOkXjrqlR16kfxf1hnOPV1ziFpU1FP13PMg8SJR
EjQUarRW8i6Dy7YnHEBdR82XsjVRTqL6K+B1e2fNc2F5r0rBCIRFYWsIzFD9nI5U09i7iRCdhxkT1Yc7amCJigpCxugqO+QkbvKEDZ0zPCV/U+gfjJulBcYFb5c9m/vk
FHD3wIJ6h+AVnHUnd+O++o4wcktXf7/F3H/gCQWhwGuQ9EJIPpxDqBIFB9hlq2MonRu+6k9KS/9uQT10PQ6gcooXWrSN+MhWs18kdnblMlmj1sFgsephsWU4r1Olndvp
aJEdXU6XXTVGwkEj76/qj7ZV+MD9MKizsdhTONHtVnNZq+uEDpWUBuzA8gfBPD92dvpwuwDiDAPA0jDqjZfJvkXGLoSgA/CfSmQ7HFWtGmoLWTqfeKzYeHmT1mT9uzJw
Uu7B73QIikzIEvN1L9W/qNwo8FNwLgmRcBOo7MPJKgKMoymjbMnCbU74rcOki16yw7BcWADXK91to3vDJMxHcvpcFJJzm9PLAQgzeg70IpCfvRMIFk0IMXf1eTGSQ/ON
UhDxWRXGtBXUkkxuljT7SEySKbn0FWfEtvrkxzaoIql6tox6npPn6JB41lj0ozK7U87LEw5ouHjxmBJ8FDHTbtrQRwHOxV0KxeCiAUZER42/J2de26VhIK0vaTi4at6R
K5RJpt7XjTJLTcekuF9od0ONFlHszTsyyd797ULzxkuh8qZe9fcW0FWDKEapoysJ3AtWH0thgEcLLqWxrOOQzCmginZEsQ1TTqRLaN51eTj3rUqOOiTSIdhTIMg5HViu
YrQbBGEIsMZyirwI42iOCHsUJQ70k7Me0Mq/eJmyjzIch6YcyG5WYSpQU98QTEW6pbPGfLtFr5czpehz+PPBbLgJ9Eja5N01bi8t5l6kn+QTmsI6TNV40HOSAtr1o3JL
soFs1cPEPKbyyQLr3YiJrMbJXwj7Sg10BPjbsMUtci5Tox7uKKy9nch7O4kKWSTDzHpdreDheYoaL+Sj1683Ys9RIG+5MiDCLZty/xK99N2UgWgWXlqLD/VXUMy90U/Y
ZtvXDjpec7Vy/XZdXckKY4mUSKaVVEto/LUYOh46wzSk1nlF3rvxSeQwlbMrefzX28MxqzDI5B5502qcsxYjXbPqzge+g22Bp+dJaQJvBsAKx5nfTZ9ni8au/H5bvlVH
VlLU12pq0LLNcrgRUrB5HJATyGrGIhRvAyxXbSXyjUHsEOuFOQ88tptiCd5NoRBwnM+psc/OK330mp2CDJqm+jWhUFMDHNVT3B22fWicu1eXIBtyVLjgcxPWVJ080Urq
Pko/h7LnmM8LH2Yopdb4nEb3qIJif+t7GOb467gelbB1hzdDo8JIkIYxe5iFpulpEYF5rX/Gezn6H+wwRxyzHY+DBkBlTxNG9I3oQKo3hIOqdfs5Q0/7giNmNeQXnsNK
VMZIC/B6PgzxQkXVBjskSlWOpGHmGtMmEZwUQf+HrX8uhIR4qAlacgyWwls8hwtlpC2WC+rken9jA5fw0Tn6eY5/KiK0dM7bf7ergetnat6frnC05QFk2PJCbRZq5ArM
gO3fSp8ahjEO9D5+nS9PPQpAO/h5MBsC7wqmrpZYLz5dNGPXf2DvK/F9Uwi07w/eCguU8lrxGBEpqU4PtGjxBokw/qxdDEAU2AhQFovrlzveuzQvOSieDkexG9zbxXJO
sGNggDkzwQdxI+VK+6oSkHFBWdoNHldpnix9AjePnTQQVFphjYvqC3dEIph9Buw44ApTmIrCL9sgmX6nMECqnn4P4SgKblRDCNTSKvnYBCt9IjgZSJIOD9xPe9s4MEMr
wxDfryCfp6AtQka2g5COOQ9jyxKpTB9/dREELQ3ApEIcQsJbYzjab5WAcCJXfUeOHlBzl586tzQeUagl27WfRjS3Sl4vSlbkGGV8RoEEtniO2F2uxUOb0rJdDaUXUuU3
wYnQfZ8FUERyWdaL3vQ3mRRGKCrOeNjM1MJb+UnCVNiFVZkI8G31ynv0DlXk/TXCn7iMK0yptYR+9W94drIaz+LREZKuir8T9aWoE1yHGNCqx+WgNCmwd1QXzFp5ZM88
jKM+UV//J45Ag8KcaKuwbVaN6Af4rKG1rosJlas2ghJtrW15AXgjmF3k8daHaiOeIMZYvFKV25YfCJZexavSA4432CgJA2Uvm0e7/ftO2T7Ncqi3rmYam7DmBmnv8csl
MivRZyRdAwv1mTp6FIx9+EdINsgmXDVfLtTmEO0wR8tG96iCYn/rexjm+Ou4HpWwmf6Y3CtA5E+TuZiQj8VugLSboSCDwmOwXM1KeVF45HAuOP6VK/szxYM/dpOnLrpu
fg/hKApuVEMI1NIq+dgEKx3umDuWtczcuBxHQlUtHAYvhL0T5yOIdbYENoB/GVUmyf1PjaDqbW+C/C/gDh8krWJu4OJ43r/pgsYnaHd3zJIWaR+4BfKIBH39aLUmg3SM
rk5mZAEfl+wMRZToSIyNcNJN+na4trZlt2oQZZMSQKLizHyzuYR6f5hgyTahMhfQnM+psc/OK330mp2CDJqm+gKuc3xHZeU/HfzdGqu7ZQ7cj9cU6l3h3+4QrqAymMsw
KaCKdkSxDVNOpEto3nV5OPetSo46JNIh2FMgyDkdWK5itBsEYQiwxnKKvAjjaI4Imc9/MKSSAGmzXhON+8CMlzwb+L4uuOgg7xv0ic+sObOls8Z8u0WvlzOl6HP488Fs
uAn0SNrk3TVuLy3mXqSf5BOawjpM1XjQc5IC2vWjcktkRXWkdNNGJOlLnv9lFr3xyZdiR0ligK8AQsrRvTLNKpl8I/9e9Zt9Pl1wtjV2HVaEE85dIrUCu1BVwLrKj9Kz
v404BFT05u3DgH/s3pY/4kZlPnIpxKaOVhj6UYuyrBcURigqznjYzNTCW/lJwlTYVwbPLcHpYrmjL/1T1wexuIbO+PLNFqEf1yUu+jk60cwuhIR4qAlacgyWwls8hwtl
pC2WC+rken9jA5fw0Tn6eY5/KiK0dM7bf7ergetnat5p/sOCBByZqJgrsB9PmG+hgO3fSp8ahjEO9D5+nS9PPduazjwhnUvFvp1+8yA//55dNGPXf2DvK/F9Uwi07w/e
CguU8lrxGBEpqU4PtGjxBkArrl35nyAx5g+9cGavkbNU7eGlTlqvqne38YpVZ9gFzZeyNVFOovor4HV7Z81zYcDZDQ8xqGInxH+IVP95cELwzVKpQhuTZeigPSc2a9Zq
yo2MgBktIR0UWvUi4hcelVVVP3mx/Ms3nQb8pcYk5E+ls8Z8u0WvlzOl6HP488FsuAn0SNrk3TVuLy3mXqSf5Fy0gx3wE/KxutzEjkYHccLM97StWrZjzAn4pq6oqalJ
L3G2GATpPhH5Ztc/2yKce/etSo46JNIh2FMgyDkdWK6AK7kLnZ2ROTSgglXdUqG1EBQDCb3Fbq+8S6ZRacH5EhitSXPhX0Vex3Nf/dhceRr4HPlhcnZbbNI8fPF4aQvr
nM+psc/OK330mp2CDJqm+jl+LuAv+dWEqq3sJFLFEdZFp0jpoBCR7RTLpXWhCuf90Pof+AYogZWJTvRIc0+TYlLuwe90CIpMyBLzdS/Vv6jdrSwaHQzO7yW6XjdQ0fsZ
2kwQRmxPwoYhunm1gm7rJYY0XPGAN+Aw2SPUJ/9fuwb6XBSSc5vTywEIM3oO9CKQV4EWm/fqtO/w1/qVCCYoGyK/Jfb5LxLBC2/MuCfIiirM97StWrZjzAn4pq6oqalJ
n9MEZH4VlXu1Yz2gVKZiD1JPXKHT2d1+8piBMgyr5Ymmp6sw2qxTuhhEgKl0hl2Z0t+GBiHPXH+wHOyMjO0M5KuG6q7/8OOx2KBWAbbfgWFVk4QFchb9OSt1jSv6DfPl
nM+psc/OK330mp2CDJqm+mcKaTUUcwQlTW7hcd5dEXcDqOkDIyv7RHxfx/5zrs56OwR0TtAXJDD0I+MksyBY339T6B+Mm6UFxgVvlz2b++Q6uprANKyFTbvMQXBT0y0y
ZcI+Br8lAckZvoL4Hv6BvGYAOrcfFNRG1LgzLoh87x5pL63+zBtpzhzvhlZGeh1UFEYoKs542MzUwlv5ScJU2J3FFVjvxWo9htQ4ZkplnmyL0360y0qrLdF3Bb9iRzne
TKSN2lnsiEhj0U3Z2T/zUaWzxny7Ra+XM6Xoc/jzwWy4CfRI2uTdNW4vLeZepJ/kEkUwFjsK8bLyVi11EuickkWnSOmgEJHtFMuldaEK5/00xMShiUDOhsIpFAifIu3r
k5fM+i5eU4qQqwYz7v4kRp7jf8BKyB1yhGBIGT7DEWA87+majo/AXVi1UX9OmVgftC6T31gJ9sOwnZVL263bJEBpF2j41gNa9O4BmkYrKp5dNGPXf2DvK/F9Uwi07w/e
MHho5MO6nwQqHMONgdxt/xT16ChVOYHS0+kRPH+caY8SPn349SuXY2OIdptoav7E+lwUknOb08sBCDN6DvQikHAlxAtAOTL1RK7J9kV+lRXxXWoMRr5NQVXjWJOxQXyf
zPe0rVq2Y8wJ+KauqKmpSTJTnrZbX416dVJZAPnPsnhST1yh09ndfvKYgTIMq+WJXMWdK4sYPPDBzpa8ThpGzNLfhgYhz1x/sBzsjIztDOTtd+qgHWwc7c+a6A8S5VpB
VZOEBXIW/TkrdY0r+g3z5ZzPqbHPzit99JqdggyapvqrAjWQ1Ex7JW46jA1yB2GuA6jpAyMr+0R8X8f+c67OejtZ6p+4BKNui3BEh6J3qMtiUffPP/RpFpYIpIxtX3Es
U3RvVhFEr3WcTsLEIUMA7K3ZDoKhplgZD7OCvx8/QU52bxpHfjTSVHLRf3I6cSxoeaxRvF9LhYy/ZKKURqMbvFJPXKHT2d1+8piBMgyr5Ymj3xXEA/WrZh3LrUjgoVBb
0t+GBiHPXH+wHOyMjO0M5KuG6q7/8OOx2KBWAbbfgWHkqUrUcUCfBxupezR4ag+svSf/byC2P+ycXnRtYAbaZs04xex6tb411BZBoYnqJLSOn8fhzF4eSjokyrUZevZV
2L1hPX3qbVCRANNsDPjKFvnuzyvnERQqz/fAmbwDVDRWY1lLh8GMnGOtxo6TUN8vYWmTLGZI6/fGsCEF6+JMGMQfjfZCWyIDqtnu0CezlMJQO6P0Ffi5bhAiJhKTLw++
SJXhkPjPkUvvd8vAYbkxb1W1RSytyEkPvyW9FRZctC75Pq7QHZZT7qBmRI9Q6iG4u2CxxrVVY/QAkeILJO2SkoKvingN87EBVSbLH7joizARgaLxaGn8OHVSHLOdrxCI
MV3DSXmD9zSEpIpSHEj8eZzidqvHNiqpzuaRkIh3gxq3b/wvYJ5i5vMaVFPIEWn1zioiWg16mApuqj3kgOdwUmIskL9N2liw4AnrfbwfW8RT23c2gkLpVz5+uOtPgmY2
Yl8EqqTTnx+JY/A7hsZkEKqaDIEn01S4utfqdfhWOLxb6U/SIUCSNL3T2f7F3nkq+e7PK+cRFCrP98CZvANUNN5b6tDFtNM/4Gd9G2x59codk9lX8HwsCw9ydEsBMx0g
Njs1j1W0KnL4BhjoV6t8mOcgQpYRuD5YllP7eHdrRhXE498u+QRSN6TYm/dEezxpLVkmdhHzezXl3gwVboahySg+vrW9xFhmrvHetGFVZI4+GJdTluLLpfCLeaVVxDxD
p650Ou2C1kIlhc1wkT221ukFPtHynGs/0n943ATy+6lmPDOskP0QWNSEXDASHQ1gxB+N9kJbIgOq2e7QJ7OUwgRA/1oY7wYSNXeAuyhtMsRDzBiIxBgukMi/+WTN+j0K
LVkmdhHzezXl3gwVboahybfp4yM5X+VTS7AahqhbMVep8Qw1FhErJP7l63KUXYpqgq+KeA3zsQFVJssfuOiLMH61d0UpAJW/49KglGZ4JxjaqSQH0rzJWmJSnR3JLNF8
bmn9+YaqLl/3K4RP/WTkqewsFtbzCrqnRjavt9F78UstuquP/W124jQlMEL5GpLw5yBClhG4PliWU/t4d2tGFRStF0Dmso/emAINisMFZVRi4vcBj0YG++JtKHtoi+CF
xB+N9kJbIgOq2e7QJ7OUwmt7jNcrLs4G3XuBOTFuU6wNbeKvLvnyZObPx5fvQFqI0kvR/55Qa3ysPeMySC/MD5qIIqkXbE3PS77K72FN3CHkAdBNcg6Y13iQjOHsYpyT
tRMcKlJDZqyWt6tbZQNkJkYP569be1iAVAHk+WTSGvOnrnQ67YLWQiWFzXCRPbbWGLKcFRFe4qFYFYzOKqRP6kbwWS4nDUYA3Orym1NNB/8NbeKvLvnyZObPx5fvQFqI
0kvR/55Qa3ysPeMySC/MDz5oQNe+n+nIgIdNOan2KXFuaf35hqouX/crhE/9ZOSp1yF04dT9+n5mrGDngPjxBE7GY4BLb6qbOWm0VRfhQFanrnQ67YLWQiWFzXCRPbbW
SnMUFLUyvM3amQNDChbP7VwuEg9V7LH4BC2X17zaFmy1wz763vulT3mf0ItXqIltuYRC72S74QhIs4oorjnSa/MU/GrLJbQqAmBXMz/d82357s8r5xEUKs/3wJm8A1Q0
Q9gdQ7+m02irW5k5bremB/nuzyvnERQqz/fAmbwDVDTeW+rQxbTTP+BnfRtsefXK0fJS6qwmHXfmjcI04SlWBw/2FvCqissy0i19HQ92B2nvam53kCcC75Y2Wf0CSVQd
Ce8tnOo9sTRXFi66jhm3HEpIF7bvNNdzxLLobrSvexUEB9t/jQ+5EraAl4BaC5mKjV2DbAwkHfg+xWR4RAyWlPweUITnVvGHIx20WaZiamN5JDuXeJ54oTkQyriWZ3kK
RBZXKnzjYNfbkKCnBaaD0nlCyu0ZyYxZcR8UbK1Unvw7d5MbdbyUWtrUqpIE0vFVkYW//v2fiN2kzX4QinWiMvKV6ZEgd6uieWwflEwQuVV8tx+BDwglboIWgaE5yV0n
BdKOF+af7KcgoK8QtnOhx/weUITnVvGHIx20WaZiamPxRJ4UvN7lyBOYsMY0WykydkprgxL3BeSu/TtJdH754+64YknRnMr3cjxsGdvmmXK6MqrstvmLGHlwb4q2xjYL
yjXiIFo5tyXfuT+wmGvR6PzyqASuJF47N6kZoEWquC66MqrstvmLGHlwb4q2xjYL9yQ2OtDhhj86IYOvjo+6zHy3H4EPCCVughaBoTnJXScYX2HjEg6snRk6QNzUJ8KN
0P7DlDXE5BmvxyVhA923cY3WUseYTOJjnm586pqEQkz+dNxSD37Vf/ohXAm47mzzVGxr/uPseIxJxHhRcT03uw7f6diZ6LcPrbzrI1dj4T08cz+tvo1nbPWPA6KDv4Ik
uP2/D/RWtMivtdrkUos87qmR7jZrxq8NryvyQpg5i72PR/X6VDIZ1AWmJqxnLiabycPURkjZuoWz2UrHkxnK89gzrj5283Y+vg/NDjPfb9RLbYTiCDt8iUfqA2gWgnQy
xNSFS8e06LGukvbC7k9C+585npdLTETumgPWcI5251eu6rySlHm+Z9UrwYJkMfIYuwOPQ25eSAg3nYe6T2QWQY1KkPBVAjB+reQ8JMujGcLGc1u5bmQ/VEoIYbIMpEfu
HLKwXL/QyCom/ryaAfo1ImaOHwTW2N3QQsWXcrFqKAkqOgZZ5jBVdcTL1UbZsjuN4hS33ZugdHKpjPuBZb3TCieDR6wbi+B2heGDRnqNBqpb7hP0Ue1PttCB7/jzNTrx
iPpEDkxbbHmjDDdZHIB6UeV8peaPFpg3KfbtF+38G8JezVetg/6x7kmRZA23GoCDyE1RjAxuq/+bkZ1mahN9IRaATFz8Bj5Pq6sT7vfisEmVRyExmtcUy8OfCy+tXIGD
gGX0KSc+UeHXB9QjixSeizrsqFiTB7anPTLYHBkpct2sYQ8bF7mxB2Uufk/jUYN+y63qLPTFasXuXIL1H0zZIHBcoxi+7YRE2ux4ptenuSpRQ3Dk70dIJMD9tmqpBYl4
ovJ2naAxmD2qiFLpD4Lv5zTawRNUd1m7rwWHtsxaifN8cSCoSBYPl2px0fshqsB3xELutIJWHTCjBxLhxlBV0GYli/ND4jvTsVaeHtwN6aJe9b+7gIPjr5/ynJ2WBCaY
hc4jSwzDsq2W8fvr8FGgKmVQmZdvpf6abBVH9k9iBBIrFM6Xob7XPZDlvZHkOHdch3w7D+O5wZpTTARIc6l7V7fLrVK+DIJehNmvfxU5rPChFCkq+kCkeZe9szRRl7BQ
VfQyYIvnWB/84gKvmFs5vshJVb59+687ImoOFPgUIA52bxpHfjTSVHLRf3I6cSxoixg7OxCB5qX2IphBl4zYXHey+1FXTJanNjZ7Wd+18y3srVjVoLBpDkXNJgjRtB4b
gJgfC521AfTaZspK62P+h2rGntEqzz6iFJTXyzRcTMB75HZ3LHH3ZzwfoWzOfBpvFPXoKFU5gdLT6RE8f5xpj7ToFjqdOytPWnzGYZTEAjAHSpB21dS6OF93vpCkF63/
FPXoKFU5gdLT6RE8f5xpj3U+e9StpFjhayEgGT3LMqZGz/J84cIY7vwp1XgSYRzs829ez1zl/6SfIOLaOfUCiPYb7f6icXS3v42NQrvfTIEHLSP8+wpviJo3VqNh029I
FPXoKFU5gdLT6RE8f5xpjxF0G9YWgG3HDpgMMHl0qGhGz/J84cIY7vwp1XgSYRzs829ez1zl/6SfIOLaOfUCiJ0aMbSWs7fsSoRqjLo+U7AiwAjNR3K7hczl6uQqYORl
829ez1zl/6SfIOLaOfUCiE604zQHFv+OLxjADjB13njM97StWrZjzAn4pq6oqalJdw9bTKh9EDRifBCH2oodkq/0O42loPNZ/6SjlCFgPKfvX0j8l14Uu+Ajc5CHf2nM
FPXoKFU5gdLT6RE8f5xpj4wUsTPFf4ydrr5XCVvar5VGz/J84cIY7vwp1XgSYRzs829ez1zl/6SfIOLaOfUCiHRUM4lRbtxL9Y8uw/z8JsQ13owzGuoiI+vUs1FIGYf+
829ez1zl/6SfIOLaOfUCiHBNDh6uLfKuyoP1PGMhe5Vqxp7RKs8+ohSU18s0XEzA44X93z6DP2CUy5i57Jvfh4YI1TwqgutfyM7mRWcHdHcLyrShRnvTy5qa6oR71dvX
4Q0ySaMouI+QcSpFglNhtiphoGPUiEgHACP+IQb0c4VOaKraJSKZwIl+/cSTgDu2cM03BpFCvK8Z26LQ1BYYk4vTfrTLSqst0XcFv2JHOd4mDtEO2m1EyFkPdRA8RgFd
hhlfr4S2FnFobWYkqqfmN6RnTXzYaZk3r5groYPMHTLyFz3rrozq9oNjHEVapTlei9N+tMtKqy3RdwW/Ykc53t7Fb4Z4twyoi3FlK3+3eMsUjZbRs3x8KyY3LFe8d0us
ek0fw4U2yAQCG2+D8uNkhfbm4Ett5WW0FjMkYuDksi01cbsTBKho0QzwH7bWK7OcMpAEL7YIQYjznEQhVLNBBgBFlhlzC/VEvIiDSHLEYnoDqOkDIyv7RHxfx/5zrs56
hcyU+9J1TdIBcr0sxXjNRhT16ChVOYHS0+kRPH+caY99vHWVYu2Pf4cT5yHCHyx8hOW/7qWplEO4aiff+4ZQVhTG/oKqCoC9WQXuTSFJ3TRrUGya8e7RAGKmFHLDaoUh
vBOy5x0+Ud09FldszMP0TsD6TRnEkLVE1gYWj1snGq8BF/z8D5v0khcVqLbanmBdHpMjGFz26BfYa8+6XnhyBeiDmjfUHWqAXZkFTZSx8trit9/poraAXU6qlNuZrHLI
f0edUXUG/8Ko7rCq3aKplhSNltGzfHwrJjcsV7x3S6xT3f7LXYSLfqJUfneAXD62qsGP1RcF2wFoZNBEWHnqrwvKtKFGe9PLmprqhHvV29e6xEH8sNu8bJ4EHOH0byCY
x0xScPizxK+Ib79tXFt2h8z3tK1atmPMCfimrqipqUn217lDJFNNYKxX6+gXOPsdVPD27DwiiVLy0qrQkDQYS71o/kjVtydLE3Fa3Ypi8qmL0360y0qrLdF3Bb9iRzne
U93+y12Ei36iVH53gFw+tpVjU3JdbypCBqA+9/rA+UMDqOkDIyv7RHxfx/5zrs56pHVOYdJ0JsO6qSkIP7hH/MDygYfjmvInAHeWWCKoJJ8X3ZYonlEbcgzirlBQ0GIG
SpWYO885l/mVBmDsOfi55V6ye5RhH/VmJK618muB3ZvpKLgzcivTUTF8EZLBbK+UC8q0oUZ708uamuqEe9Xb19zuuuA5XKeLlTcnkr7vlXk+mIQSFz1raxKu0b9je8vH
S+MNl5+cCTlYD98T1E+4fr681kU0hPR4xNrVFy3ivRnCFAButZaZudXBl5oTDolOV/fMcU9SrRlu5ZGKFAx4CK/27H6GjBWsqsrnykHeIMcZgxfsCYA7U5Vc7wXVUfrk
VAKX7ebETX/uQIIcYPI3SUticIHi89ORE55Qc13XAyyvzyyV1naTFDy4/PKpNWOhBbTucZXm0vmCp+tI/pUK3JrDFb529zF0DOWTyBydS/hjKv5MjCl39bl7OFPfi+0+
xJof7l5jCI8AxY5paCL5GWajUoAjIAdZlPH2JS61AdjDs9oyqeCLyk8heTP7vAWNkNKZwWPvVUaHSi6H119ivzezRHly6aXR0kHKfCP2m6FVgPiY2yMqSF5Erg5YQYMx
/4y3qGR66K53g9ijNlcMI2eKyDT29qDlDisDyetq+r8XA/9Wj1rav7x2Mv1I7eioyGfNfmYuskyU1LRQ4MpV3Vf3zHFPUq0ZbuWRihQMeAjBpXE0isrLAq3HbN1BIxWK
9C12vCkfFDZsDcjRw7/Psb0mP2daVcH/sMESlhbvFpl6qemdLkQkti7F1xCmWuw1oy38hR6FOJ/K4D9HrDtz5/yKdveJmrnGYYsQ2nXAuu9is542Vyxn1qQ7SX8LKIcH
zWf6gYMAm6EsDaoleE2RQAEISxbamfK+Y0hFjHZx7Z2+CGgvGYTEhE2TRAn0aMVPShjtxooKbwNQkVXallu07YssVXNHx1HZ63DqDk9ZOnDsvI+shJYKWTuUjBKQ4cJA
4aKagJ2SbTxSEy05sdDQ9n4mixzJhAoJFVdHKqnmK575tFB32Bth6GfX7kOdhpUCavbzzhXRU2TtdBLsDjCxqIROtuN6mcGxtOTbKtXiIjhX98xxT1KtGW7lkYoUDHgI
RtMVBk05YVXveZD+zjFgBTaX5C4pntXfF/xP7IOlB87A3ggbsFtxbvAe2lFvD1g1LQyfJTyKVp3fEBmHHAHPsOZNT8wVJBWtszyPmdr5cyMkFOFESOV2J4l76FonmJ1A
AqmrE+knpVw/pa2cGiLYRS2s7dvKXohNslyaEhodgL5vkDEK4WfzyV6Iz0bTBJPmO4Wpjx4o9qxP2di3afoCWDIr0WckXQML9Zk6ehSMffiNcu/MvWVC6g8goadN6PCQ
n3TWcJ539LkyWOXIf4O8B8D6TRnEkLVE1gYWj1snGq+XUAGBuXiREdqmDapXBvT6eHXB8bDFa4ORkjIjwyY8rC2KUpGiqla3dh7es4K6FishOiqx6HdYRXlh//0c55dZ
GkF1KwPBjmA5hmyqmw2zfs49XXOIWlTUU/Xc8yDxIlHLqgBaqXbq2pPIUIP4OTrsXY+CQpQrfyd2QAWqA6ZEavSeLK8+NBKsn6wDYLTx0j1F1vwL3t5ZaytTrASaCQlr
HauMVnT9LaYC4ImXaJuH6rH145SDO8LUillmLUv4UOqdMoCRqijYENYbn4+Gvzk2ZqzRoERlCh3J4ktIQWU16JcgG3JUuOBzE9ZUnTzRSuoGuqpUheFQ8+zYiq95hzFS
6oZi9vUPZwN5tH4jR6MsOXeuGPCz9k08GICwMQGrf6Q5wkrjf0vOptUF9MN28RBUJPT4itwGWs81NtMkI6CapQ7nnZHUX/zNIjBLAmmWcFgNpvvSzSF5rkx8LZA97057
5wOsNlKACTBp6rPhQmpQWzDDX6rfRTIjs9ijnhoeKaOwsdvLGXEhX5S8/XjhK9U6UpEQgVwiiiqeLFIDDOKg6lT2MHUVJ9f7D9XBsP9EI+mh5+Nk/l5icYZwUUyYYUHn
PIk6St3x8Wvl0Wak0EvI/2MeEfdrNFGJP+V9wJNVSYIiFt6xH84g3MSJrvrCPYQe1q6+KAwHSgBPtjS7Wi9ItAlxOkkDM4O5vSB73u1RwQTK2/nnO6BNdw4ME6GofC5C
qygO3i91uzT83odDQ5ZjYCsUzpehvtc9kOW9keQ4d1y0LpPfWAn2w7CdlUvbrdsk6USS1Lj2YD407zf3uRMbMWnn9A6AjFQUyXDeJ5M2rNZ3ydDPG4SRxOccVhtsdoaR
GUDV4MNdtPwwpbLZTO3kqxh959RFLh8eeEaDVcGtMP7GeLwmweWs3oQE37sjYcCiVj6DoRELoLb5UrhdXmYj917YCW+5U0zWocD0f+cC5c1pY97WvnTF5W76zFz0yS3S
FxSguGB6vdKi0ltPnUiETovTfrTLSqst0XcFv2JHOd6s3qnRGnxdsbU81ZgPbrtkExfUgoJ9M6QCCD4czwcEmLuwqqT0nDjvfGzptzrFz4uXTQpz6ISLdQs7f6+95C2v
2PkBGYavwQZGWvKnKuotQhT16ChVOYHS0+kRPH+caY9+LO4bz1CxAok4dfQTV7YkARzvl6CkVE28hhVpwzTu9YTlv+6lqZRDuGon3/uGUFY9R8HcClQE7hWaNXkIwhYP
9k5zS4A8DkOAJPo2ItdzvgOo6QMjK/tEfF/H/nOuznrfhrpInfvmA2WKey3W8XZaFeIPMFfmw/IE7XO7oFaibwvKtKFGe9PLmprqhHvV29eSv5jIdVqwbnNWKxptbtSg
ogQ93u9KOIesbAvIGclFOwvKtKFGe9PLmprqhHvV29ccseELrHcUeVrfGCcQFpnYyOOkWfDOHs/YKl70hVnudQvKtKFGe9PLmprqhHvV29fpjom7a3hS0ZoWybojsFK1
4XLS4kIeLi5AezlfrPiZ0jDNOswLA9rSdRp+HZAEsDZ5uVQa1JAWDrpuoGCMZou12QoaTnPwPuM/8ePEiEev2LiqtBkNzBa6MNy7BH4VShV5uVQa1JAWDrpuoGCMZou1
w8uYYC1gFLHeba5z5/P9sTLmR2YA3WXL+4qN2jWXgPzrtlQ0hrlkhrjul0zdsJZ3aQf8r/oexc00rJzeJCScg7FN3/4OJZktx3zb4X44rmd9Vfz6oH71BpUsazyAhgrK
0MSPzr3MXmswE6n9jmqm0/Msm6nfH/Zn7GN3LKatcQTcRWtkbkE2Id3ImEB7qTqtXyhCx+9A62kvqfRNOA2IaYPOX2eJT9Jy0C0NflwOqPSxiHBXLgkPh/UDjMQSKXSy
nImU1ca24ri9Pxh4pMs5eNIkTxechcU/PykN36YGSMxC32ZSD+RzzCNuAIBN9Sjvf1PoH4ybpQXGBW+XPZv75CgkX/PrQYSxk8IH9U2/t3mbM7W2Xv0L2PQhG3IcK5Lj
LCuoG72kJ5yEGoCM8L1GkRB6p+wDkolr1psQq768M0fndMZZfWDbhyOZPbaja/Kl3iX5Soaiu0TTNS7wVkKcqgZU43IzZbAzpjWmHCSHPpBqxp7RKs8+ohSU18s0XEzA
OlESjkwzCV8G46hj7zPQv8R17SpVGWcicFtpHBHUYjFXvrZpiPDmOSJ8tlM+R4UXbJ8rT/IyQaRj1D3WOHJrxCkBZR8Lb9hIlIVtDdztv8LO4R7MEu6LwLgXj7G6y+ft
1kDeTQSet2EUifMY1sn83J+onRTU43MhnRaHMYxZTbIlIgE9YV7mBazsxDh+U0/VhCYQ0A3GL17vDt7+JwHti3XAuhRiOcAASPBoIGAJnoo1zGybZgZbqC1AxRURnjP0
B8W23qMGZmv8OFWspkInHWdyQjWL9s7MOjuGNxYddac5kg5oBNXlZpnT78BR9Jr6OBp778zqdx4K8ZUMaBg/fT0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4
Nz0urYhhHX+R4ghqGOl1KD0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4EKWnp1Qr/3FaY1/P8ykJaF41Ohg/0LmMlfcE1HmZfCqRpQjoF0MHhwFqQCq8NNbS
ys5+d1LWLIUzk8A4UjJClBSPLhT5Ug+zYUNxPYvJfBCrpY9OqzrTG3VR9UcCk3LYnreOuqgKTuhm8gA8sOhYIXyEIcONU6WLfxNRUuK3dEZ9UnWNv+qXe9NKNetqKiML
h1mVRTdQuGXbKqXcRIbxHKxPMPwdHZ98fQd0hkImXYy5FADXSdbwZyzUnjosLYDgtpzsxfRgVAH0LvQCU/Sx12j9cy7XxalrE4vLfskOs3r9WuSPBxbbRLmWDUpcD6+K
+ieDMgKtUjftuTFfyYFyqWdyQjWL9s7MOjuGNxYddaehHAwaaptY5hqQTlsIrzlyyijZh8LmwfiKibX/WkCyZDRi6/Q7+mjbCiqWtUGmNqwnpct/UjXD7BYTEByjkLBm
WUL/mIf+SHBl9LwlITGIHoQmENANxi9e7w7e/icB7Yt1wLoUYjnAAEjwaCBgCZ6KMNTmHVsUf/ipnKBod8eu3A29QjKh5tOiuQYB0wXkQkN9RShOX4pAd5/GmofNusGv
8WYCQOe3HM2U7TOn57FjPJO3R7iiZBl66Ipf3I1/X7Ud+F915PH1o2o+2tddj/r8DmlC5SuGORuXNB46ezok/kFZlrk5Wn5ffewryhLrNHAHM/wMyJggiL17wuNW4mo7
dcC6FGI5wABI8GggYAmeigEFWBYWc6Ue1zxHl6BbIVWIElWnRABGIcVRuxhCs124q6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCEPnNzzzIRNI/WmkdpldLcs
4cxe+W8T1i50iFuqTkMY0P9aPE9sH7MI42fPI4d1a3m/bUOMp9282Mxd3WcLOGjnehl7fm8lNETZlrm8G0tCIf+q5nY7WBv2SyrLHBK7AUhI1mh1FNCh8htDhUnJ/pgZ
49FOnDBDSKeL7UkwD6rzd9IGiqxNdkF8pLgKpY2b/XsGhtgRD42HToRY059LAeJjP+yrZrzb30ky5gr5Y7KjmiS9jmDHu1Qfdsy2GoPFOL7WQN5NBJ63YRSJ8xjWyfzc
WDRRqamA3OL7tIxhV/DqUx4xXI31Vr4NLsGmYO2rXFi2nOzF9GBUAfQu9AJT9LHXaP1zLtfFqWsTi8t+yQ6zeiHizuNfVt0XxAh0L15EPZRY9wCznmWd6+J+VM72M9b1
fUUoTl+KQHefxpqHzbrBr9lhXiI/K/GAWlHmKT5vFxlptieiqqLJ4tCYKHX6Rno0UMgCsOdd3THJRr23GJArZ3peWNBb/DtnXcivBtwoaWcQD7v5N9prmdevrLW78W/S
Lhbj3zk6WyHhfzi5rOaeXeL8ZcPWLipLxcAp34JV9fYOaULlK4Y5G5c0Hjp7OiT+dXNZyUTTzsJbpasyc6kY3myXLVfUsrBS82yf6HR7P4dl5WrIRc/wmYmoQ0+8L0gy
Z3JCNYv2zsw6O4Y3Fh11pzmSDmgE1eVmmdPvwFH0mvrHd2cmkEXyK5OnbigBhpLezuEezBLui8C4F4+xusvn7dZA3k0EnrdhFInzGNbJ/NyfqJ0U1ONzIZ0WhzGMWU2y
Sovp5v1Q/Ic8eGjSVSHx5OCn7fFodktlECJvZVCGvc+2nOzF9GBUAfQu9AJT9LHXaP1zLtfFqWsTi8t+yQ6zes4zLCah9DO4zlitHEIUDbbOSfxJs5KIjnFm9wpryP/A
kaUI6BdDB4cBakAqvDTW0srOfndS1iyFM5PAOFIyQpQ6mHABMu1oDkLQSgigrVX0sgtCseZlGb+p0hvkmsHk4R34X3Xk8fWjaj7a112P+vwOaULlK4Y5G5c0Hjp7OiT+
M6Z2gB/d5bO4DGWjQyfri3IWe+hWVaroxeH3J+FAhSsNvUIyoebTorkGAdMF5EJDfUUoTl+KQHefxpqHzbrBr/FmAkDntxzNlO0zp+exYzz1FxzbbSosGnjOU+7RFFRf
fVJ1jb/ql3vTSjXraiojC4dZlUU3ULhl2yql3ESG8Rz/w4vxX/mfRPtiUY9y2S8asvCxXFzA1OPPDRZ1Z+h1cPkP22nr8fJFV6efCxjqhpyRpQjoF0MHhwFqQCq8NNbS
ys5+d1LWLIUzk8A4UjJClDqYcAEy7WgOQtBKCKCtVfSpOT4FnZPkKM9xG883Se+Oq6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCHTurt2nFZaAkRvFI7la4G3
G0R/0ijoi9s/fJAkXjJeT+HMXvlvE9YudIhbqk5DGND/WjxPbB+zCONnzyOHdWt5v21DjKfdvNjMXd1nCzho5xACllXrM8Iqg0kzbxBcCdGogzoA0JCEC9LEOpoGM2L0
NGLr9Dv6aNsKKpa1QaY2rCely39SNcPsFhMQHKOQsGajA53GfIZT5smblfKSHUslnUy/rw9s0f4sAG7ricWykpGlCOgXQweHAWpAKrw01tLKzn53UtYshTOTwDhSMkKU
OphwATLtaA5C0EoIoK1V9I6Cu+UBSm+HeJxZ6s7JOxCrpY9OqzrTG3VR9UcCk3LYnreOuqgKTuhm8gA8sOhYIdO6u3acVloCRG8UjuVrgbebawVLOF4aRPvfBD/rIBNJ
4cxe+W8T1i50iFuqTkMY0P9aPE9sH7MI42fPI4d1a3m/bUOMp9282Mxd3WcLOGjnqi0pg/zmrK01iu3SyNZm3bPmkhWtsshVg4hEsAzRVqk0Yuv0O/po2woqlrVBpjas
J6XLf1I1w+wWExAco5CwZiNjJjdqUXse5bxrRXANiV4pOsKjCzPm1ewlFzbQjbrlkaUI6BdDB4cBakAqvDTW0srOfndS1iyFM5PAOFIyQpQ6mHABMu1oDkLQSgigrVX0
oXu1jwrYxABC0fgZ1/Ndlj0wjltC+rQNEVP1Kn/fNi5pjdJ5wfPZn7ICmeoi4QT4JyIU0B8hrSosy+pP6V50W0WU4NvZCUUdqIEukdpYb32veyi0N13qZ4pHIXwmOETs
el5Y0Fv8O2ddyK8G3ChpZ0B7/I2uW8yCAgd0gntygkKfTMTkQZJtmqystSAJju9poFrLK1cGWGvTwmgQHRgnl/3DkbC/vp3zYTAKcp47CuNcMiGcHLlMTCHxO18O/hmm
C1tl/NHhUsKnZWwQl8ghBsoo2YfC5sH4iom1/1pAsmQ0Yuv0O/po2woqlrVBpjasJ6XLf1I1w+wWExAco5CwZqikO8XQ8Bb78lzeeDnZQ8vR6QrQKXKuHihhWoz30oUV
/6rmdjtYG/ZLKsscErsBSEjWaHUU0KHyG0OFScn+mBm8gCZW2ghDXdsYo4PGkYs6q2npqZswr7PCz2avnGW6o+Gk+cpWRZ0+HogGFpfVNpg0Yuv0O/po2woqlrVBpjas
J6XLf1I1w+wWExAco5CwZmXqmdBZ7MbNI829S7+XXf8uFuPfOTpbIeF/OLms5p5d4vxlw9YuKkvFwCnfglX19g5pQuUrhjkblzQeOns6JP51c1nJRNPOwlulqzJzqRje
IrSdQm+FrShaVenAAMyR3psS+RSxFHong+icBPGETZuHWZVFN1C4ZdsqpdxEhvEc/8OL8V/5n0T7YlGPctkvGsNOGTQdJtu7L9K4mRCRvGkcfDHRog9fn3kEy6yNbSQH
0gaKrE12QXykuAqljZv9ewaG2BEPjYdOhFjTn0sB4mNSTRej+I45HK0oqC+8rtFugfwF9bfsmVjLtc/IA9l/LoQmENANxi9e7w7e/icB7Yt1wLoUYjnAAEjwaCBgCZ6K
AQVYFhZzpR7XPEeXoFshVeOmLbYtQ1xwQxA8pELFrEQHxbbeowZma/w4VaymQicdZ3JCNYv2zsw6O4Y3Fh11pzmSDmgE1eVmmdPvwFH0mvqjfsWuKq5lr+IihlDWJbcy
S1KFdSPx3E+UcDsogbWtuKulj06rOtMbdVH1RwKTctiet466qApO6GbyADyw6FghasivPMhniWIZoZ18kfiE0W6D08Lj6qGAapn5oZHpJScHxbbeowZma/w4VaymQicd
Z3JCNYv2zsw6O4Y3Fh11pzmSDmgE1eVmmdPvwFH0mvqjfsWuKq5lr+IihlDWJbcyEZMwMTq7cSnoAad6ZWG8t/+q5nY7WBv2SyrLHBK7AUhI1mh1FNCh8htDhUnJ/pgZ
suGgY4ulq2aX2YKDLM1hI9gvAFKLs6TojOzjxO+UUtirpY9OqzrTG3VR9UcCk3LYnreOuqgKTuhm8gA8sOhYIWrIrzzIZ4liGaGdfJH4hNGNGa9fO6d6G0QgnRcpiWxK
LFTUtEI9HpEMuCXZQVivsjRi6/Q7+mjbCiqWtUGmNqwnpct/UjXD7BYTEByjkLBm8kTSW8vicx9dhVihIYXbhVSxgZdCn07FuGJOJvkyAHmRpQjoF0MHhwFqQCq8NNbS
ys5+d1LWLIUzk8A4UjJClDqYcAEy7WgOQtBKCKCtVfQqd4czmmWM9eNRQz9cRjGqoFrLK1cGWGvTwmgQHRgnl/3DkbC/vp3zYTAKcp47CuNcMiGcHLlMTCHxO18O/hmm
Kb84bKX8lOjN8shLDy+EFlD7XmPnSRI3V0JtnjqhPICHWZVFN1C4ZdsqpdxEhvEc/8OL8V/5n0T7YlGPctkvGsNOGTQdJtu7L9K4mRCRvGlbdzH4i6gvrP6SZEhHe3IK
HfhfdeTx9aNqPtrXXY/6/A5pQuUrhjkblzQeOns6JP51c1nJRNPOwlulqzJzqRjeFZk7/MuNN1zKoAbvJfwbMwfFtt6jBmZr/DhVrKZCJx1nckI1i/bOzDo7hjcWHXWn
OZIOaATV5WaZ0+/AUfSa+qN+xa4qrmWv4iKGUNYltzIC7JEyIPH5O5qYtxS17R9UPTCOW0L6tA0RU/Uqf982LmmN0nnB89mfsgKZ6iLhBPhm6a8p7V+x8Cx6PT4SldF+
ZW+kV6/nv9SQ6QnqTC5n4Acz/AzImCCIvXvC41biajt1wLoUYjnAAEjwaCBgCZ6KAQVYFhZzpR7XPEeXoFshVXJJDzBfrqh69AlUJKB4+WkyAX0dQ6YECa+BLZXOU0sR
tpzsxfRgVAH0LvQCU/Sx12j9cy7XxalrE4vLfskOs3pAt9w3BZXKqVM8UkrHqlw549FOnDBDSKeL7UkwD6rzd9IGiqxNdkF8pLgKpY2b/XsGhtgRD42HToRY059LAeJj
Uk0Xo/iOORytKKgvvK7Rbij391tiKF1C7LC2pjAOIN9AK6Pyy6bZn4QdhYbHG70YZ3JCNYv2zsw6O4Y3Fh11pzmSDmgE1eVmmdPvwFH0mvqwuHAaTmMwzV7u9YCcLZe3
UPteY+dJEjdXQm2eOqE8gIdZlUU3ULhl2yql3ESG8Rz/w4vxX/mfRPtiUY9y2S8aw04ZNB0m27sv0riZEJG8aTOblJqw6+IDrzFC3yjXGXc3G856ksnOHJTvi75tG/dk
/1o8T2wfswjjZ88jh3Vreb9tQ4yn3bzYzF3dZws4aOd7WIIkQVa8yVKZoYOZ2sl5mt6PnBe86/4qmkAwLM+jNWAyZBz7me2TgqHj3Rd/Q49w/oQvDTwp+/5xsnrQnPGk
/cORsL++nfNhMApynjsK4/tAKbf6NTZpp6XVDJpbD+QSzEW/W1OgYo7nIglzb/G10gaKrE12QXykuAqljZv9e8Cd3b84K5sCXKusIxcsYqpHxyKMXvV6rkhL3+bdBcl8
0gaKrE12QXykuAqljZv9e8Cd3b84K5sCXKusIxcsYqo+9hZua3PAvG3m+BI2xEluZe1+tkcOH+hd5TWR5KBYgX1FKE5fikB3n8aah826wa8uXQphG0yHehcEETuZ/D9i
Db1CMqHm06K5BgHTBeRCQ31FKE5fikB3n8aah826wa/D7bkaZSjg31gI9RJjLKxUru24ta7dKOH3JMqAXsROgqulj06rOtMbdVH1RwKTctiet466qApO6GbyADyw6Fgh
Zlaupsu8MG6wOn0jmC39F+JSzQiRFDjRgkXAWFRr9059RShOX4pAd5/GmofNusGvw+25GmUo4N9YCPUSYyysVKHONKQ2w1hDBYZEOX8AuNkHxbbeowZma/w4VaymQicd
Z3JCNYv2zsw6O4Y3Fh11p9mDwahrX1uZJPbVEPWg1FQip4tmTuvt65r3ZpdTkk7Gz4/FGgxvRWJAkqCorzraUTRi6/Q7+mjbCiqWtUGmNqz+4cAuvSY/V58BDExZGMNs
Gc78T2VN0uN/SWXgOLBon87hHswS7ovAuBePsbrL5+3WQN5NBJ63YRSJ8xjWyfzcBQf50QtttJhDTIeozgwvIPUXHNttKiwaeM5T7tEUVF+qKADBqzbj64TC9MYGGQtU
tpzsxfRgVAH0LvQCU/Sx11jPGARlgPg/3/jJcVUEG07QVlrKdl7zll0Z4OjusL/D8zi2QoCa5l0lJITockQYGJGlCOgXQweHAWpAKrw01tJxxs+xTuDuxt+O/bftiJxY
w04ZNB0m27sv0riZEJG8aSBhoe/FaHDGtmVg82AtXfHSBoqsTXZBfKS4CqWNm/17wJ3dvzgrmwJcq6wjFyxiqnEHFErppmd2Lz2lv+fbEYjiIrS2RcXSoXmnz55Bk2mq
8zB4hDMjihleP2SOQNKoO2dyQjWL9s7MOjuGNxYddafZg8Goa19bmST21RD1oNRUYWym/khygRnTyDM9IrX+b3t36/8Bx1DeylFB+WZpmC7SBoqsTXZBfKS4CqWNm/17
wJ3dvzgrmwJcq6wjFyxiqjqYcAEy7WgOQtBKCKCtVfQ9fE+NNh5xyPqXrsyxFQwNhCYQ0A3GL17vDt7+JwHti3XAuhRiOcAASPBoIGAJnoqha9Kx5GFHKo0CaS2Gkn39
4x0ohNxLS6b2GK/6gzx1hAfFtt6jBmZr/DhVrKZCJx1nckI1i/bOzDo7hjcWHXWn2YPBqGtfW5kk9tUQ9aDUVHJJDzBfrqh69AlUJKB4+Wn4wKZucswBHhVsEz8CH3ja
kaUI6BdDB4cBakAqvDTW0nHGz7FO4O7G3479t+2InFjDThk0HSbbuy/SuJkQkbxpiEJgifNmqqiMr28LnKseStIGiqxNdkF8pLgKpY2b/XvAnd2/OCubAlyrrCMXLGKq
OphwATLtaA5C0EoIoK1V9DozMCoodU/Zmp+XKhn1g0SEJhDQDcYvXu8O3v4nAe2LdcC6FGI5wABI8GggYAmeiqFr0rHkYUcqjQJpLYaSff20nECt8/BM/rW+28/ef3SH
DUd6urK+i4RTqLzpV5ovJnB0eGiULrs4nn6hahbR2nJ8QRVMIQ8kC3djBy/HzmKTJ4ya6GjRfMziR3ZtXVQ2iXbxmEMZX+f870ka4yabJVOorqXdKFuVZY0h1osc8y5S
figZfWFG3QGJ6LBbjGfW+8Sw1K3J53qwMkrL/BIlwG+cS0zKiohbbdnA46KuXpTkLqy/dEiQyU8H+96Sm2Kp5Ag5R28Z3CCX4uQclfmVx/8afdVGIaj+PvKEyZVb4FiE
eV0nPbIM/WRxqg5st8/E/QTi97qxVkxmLkTtQVyGOWC0t20pfGoquWW+SPmiN9yLoc40pDbDWEMFhkQ5fwC42cSw1K3J53qwMkrL/BIlwG+cS0zKiohbbdnA46KuXpTk
9Rcc220qLBp4zlPu0RRUXznpl3dsYASDkIoQ//RLKNPeI6pQYCAVexktj68ueMtNubtXJ1bOTHxT78MOolaveey1mL39dqiHMCFbE50MXRSe7j1ugJyVc2hfe6Dgaw85
OphwATLtaA5C0EoIoK1V9J1gOoyi4GCLsUE5eTueqihNCCm6LWRKQPT1MyUfei2D4nfTTrUsYVpC5EpbxrdnDcTxmSF9Ia53R93eIHrWVIm+mM0b4r0Yxl8ghQ/ZfT9n
Dg+/YG6p7pDeQXRSKFf/N1vUDIV1r1w7VPkVjeR9vWKWAyd1M4Gsj+Iqz4J6ikeKkEpHDAY00AkGAgiaeiy8Sqiupd0oW5VljSHWixzzLlJK6qUuLnBu3IzHw1hK3IFk
TQgpui1kSkD09TMlH3otg7KHEzIibU+kJhQpUoJXZXW41renR+iN4qClPsCFMOwTK4/B0ZjHlFHxaKbw7v2ye+y1mL39dqiHMCFbE50MXRQiLmTRLzhXplLyo4Bcw3lV
6wkvR5o8ExS6KbCLGkUJXvJnH9Lb+MgoTgYwAbk7i/uEmjDbI2cFpwvrz7glqxzVUPteY+dJEjdXQm2eOqE8gPYMB4eoIzzJRqgh1PAlExFlfCgWtqSZaRfowshrkHNR
DAW98QdXDI/BvpSoqVMoQcxzYWNR7Snt6cJ+Ar6MAetFRWnh1wD9jR92gNnkOnr2TQgpui1kSkD09TMlH3otg9kMmFPSAH+xnJkgwY/rMbwuFuPfOTpbIeF/OLms5p5d
k1GZnOhYwRLz80fb7o3aGvbPKFu79N3Zmmsp3seNYA6BZ7V4hIhsaVJMXtqdBoUc7YXb+MDXrLGm0/LzTX6X7q7sFiZbfPhgZz4WiRR+3ru61fu+a/dg4WITWc4Ll57m
j+iU4k+9jCY27Quh3Sdy2iIuZNEvOFemUvKjgFzDeVU6mHABMu1oDkLQSgigrVX0Ae5V9EYH/6Rct67fwhUICB1xVGgXXD6hV7BK1EQpA4xIUhBkMvRReXH03cQwv7hT
XlvMVGYbzB+z5LPE/iD6K00IKbotZEpA9PUzJR96LYN4nUtQUsjmhZIrnd3MQOXA1QotJShNGedyyvsWEWXwQbRQhLhWooX2/XH4TuGlSjlB3YGyvsz9etMepEm0ost1
m2nwJA/154b4PBfJ3YJ3Wc7hHswS7ovAuBePsbrL5+0lI6qYd+rj/TWvy4kIMMBHw04ZNB0m27sv0riZEJG8aSBhoe/FaHDGtmVg82AtXfEdcVRoF1w+oVewStREKQOM
SFIQZDL0UXlx9N3EML+4UwvUj/um+Gtb3brK+YoTUuuZ9uGqJ75QO8vCVT4pCl5nKKDL9W8h/qWxTQJnRRrV1USuqtFaC4ssy+ITOZpmGMeZi0ngoHyZlZj68oc0s+ur
KD6+tb3EWGau8d60YVVkjrtL1xweuMrDBKpLe1CaRpeG0j9W7wwlpjCqFvhZkCwU37TEmCB5IFaHGAgrYdF/GFD7XmPnSRI3V0JtnjqhPIBDDeD0j3FDeVGlN1qtpata
8iRjvq0o0ZdwHrs6rDRshSSRZ3A3MHMDQO3FXgmmEs/NJT5IBwBeGJVTqyT3XFWuwE5wpFI2s9yjVgXmnA/BX34Eqt+JrMdskB7OBx95lI9VIefREUutdM++DyhXD0Iq
HzquMqRvyeCEoClNeFN5DKu3dUBInu0gQUvkuP2C6FGu6VyfN0blWnTIM6e3PwBpSW9NF6CKBuHLdrfZ8dEq9ryXXHZzsBb4uHLOBxk5GGUUjy4U+VIPs2FDcT2LyXwQ
U6bgO2hzpVM70iDAxRsbW8DI4k6l/Kxkpzgccw97EH+STKcYjofvHyr6qf2GdtEn1GX2vT8rTyR4SJ23565RSYbSP1bvDCWmMKoW+FmQLBRIEfkO48FLi3L5x6x2N+q6
zuEezBLui8C4F4+xusvn7YbSP1bvDCWmMKoW+FmQLBTSbgqj61H/KXBe40jWoc+xlcqqjdjwSWoWWbNRs1rTYhs1ANiXyN3o+yy4EPvlPCq/lQs6W3xAGhV+3WI/bZhm
BGcD6shfv43FTeAoRSGd4GLw8EONRTiCKVwTP1lZJpXFi5iCRQI1fX9c8gM7hiRGkYWK5rhg4F84Rp6yiwhWW9VEJBF37SY2UkbGUp6lns9ErqrRWguLLMviEzmaZhjH
mYtJ4KB8mZWY+vKHNLPrqzVL+8pTMAnPFVolZIz9PIJVIefREUutdM++DyhXD0IqHzquMqRvyeCEoClNeFN5DKu3dUBInu0gQUvkuP2C6FGGafkjOWEHww7GIaE4BWaC
wApdfrcKTv6PuTHpfHsrHbZ2hK30QwSc5RdYQQJiciald2okJwSCqX7JfX6XQaVCBM+zh+zUAfEtGxg+YznVe0e1Z99X9r+dAMMtGfkok5Q8FHHoPOMEX0rapVgM7ekH
j0de5McOYi7kBiq5nCP2wY4R8zJhe3kc+ZAXe6nIBLaYzO2NMW9cUGcfSSwE5Az3zuEezBLui8C4F4+xusvn7YbSP1bvDCWmMKoW+FmQLBTSbgqj61H/KXBe40jWoc+x
PedopCWnyGgXuRkNXmWpfM0lPkgHAF4YlVOrJPdcVa7ATnCkUjaz3KNWBeacD8Ff21waa0ncWkDBYc1bolwruio0kjYRofXmlqdnWqJ/5wnATnCkUjaz3KNWBeacD8Ff
bKgTGeSCfbr8Kun5OSSfk1AeQeaIM0/FlxZ/+B/DSTsEz7OH7NQB8S0bGD5jOdV7y81XMastZPEN+1od/wQUjUHI7MAGWbxubMxfE5k58NNJb00XoIoG4ct2t9nx0Sr2
vJdcdnOwFvi4cs4HGTkYZf2t33p7MFwsnJaYWj1zdq/k2fuhZJ1Od0on+GVgtYnof+GmioSgrNlSuaPcAG0tMGEFf4YMd0AINRfh2BapoNhptieiqqLJ4tCYKHX6Rno0
qXrofZU3cRW/vOetq21gIsj+T5P8di6XieeA1YJl3fqOEfMyYXt5HPmQF3upyAS2GjiCMGxE+Jhb43u6l6y29dd+FmzdnozwrEFseokVkY9ErqrRWguLLMviEzmaZhjH
il611u1RgfZ3Zx42nEM8bEfHIoxe9XquSEvf5t0FyXznIgz052WWswq9py7tYm8LiTcIMIvt6DakCbSACrs1xshaFgYkKUfCox9efB7JF4caXtZ2NI2+vSnggS77H+e4
bR0ky6XrOB4czEonuEuRisCCJ40EwuzMvswHajHVVpAEAryO2LIZOMoPRLzF2cA73SqR9IuGx/LgCWP6V834ydbwlwLwkjjSm6zuFCtbAWVjbSlVOvqIF4DXPbPPo7rG
SW9NF6CKBuHLdrfZ8dEq9iOSny1dyJuioyGyf6XXcLX08m3naMyF5bbVr07FQEGzycV6tcHflEWqV44XHkGI+b+VCzpbfEAaFX7dYj9tmGbhSVQdq3JObGBOxbRH/cjC
5YulsJuxllqZGn0v6sEgA1Uh59ERS610z74PKFcPQiofOq4ypG/J4ISgKU14U3kMUk0Xo/iOORytKKgvvK7Rbh2i/wE4d0j+T/V/aSo1cQLNJT5IBwBeGJVTqyT3XFWu
wE5wpFI2s9yjVgXmnA/BXyhsExIsXhv5uooAECPCcEUQ/x315mcsgvCl7nQpaKtEKjSSNhGh9eaWp2daon/nCcBOcKRSNrPco1YF5pwPwV/nni2uiPG03BOTqTDCBQot
CamxY8v0vG9RxltMISRnyBs1ANiXyN3o+yy4EPvlPCq/lQs6W3xAGhV+3WI/bZhmunvKRIkwi/kraVNWubdlpniW4BG3yxO9Uhz3CV57SZ9LNYsurzwS5IIyc1uTOM5x
v5ULOlt8QBoVft1iP22YZkXn4NfdV6FGZpAyw6JElIcaEqmnEIkO4cBotuVx6LAM68kEo/oBm0wcwdiWSKOUhcWLmIJFAjV9f1zyAzuGJEYW3hypigqmcStUxzv/20/t
1nVOaIW/xjOCitIsevM9er6YzRvivRjGXyCFD9l9P2cwas+xevyW95wK+JCBNMp6VSHn0RFLrXTPvg8oVw9CKi5xylCSuvwyI4MWq3mB+s8HcFl4dxQKD8838hggYsYC
ggLOmCPkFgXqsyNh1JZ0hY64hFGigmzSxv33v/XbSZWdO7lPv2l1g7sUl+EYXV4bKjSSNhGh9eaWp2daon/nCT63cZp3PqXg0oGwM/iY0KQ6OgLsKZXP2ag3lR+wLDyx
gKQMd1BdoggKzx68v8CGK1MGaha5nLTIlr6IZcRBn0XGL4Lvq5kYFRPTI+U67ChzRK6q0VoLiyzL4hM5mmYYx7+XueWv+aVxqYz7x5bYBR4jj/BKhTa47wYhUkLt6bsd
68kEo/oBm0wcwdiWSKOUhWx74GoJyO9XEjmz77yLuOF/GaAOYA+ZwEi8nCdQiBA2U6bgO2hzpVM70iDAxRsbW1EDGRwjfzqEqzhjMh8hEa2h7o+mpVU7/YTXNBxL49ki
eMVAb5PIGZcO3K9bguJ2P1MGaha5nLTIlr6IZcRBn0V3PgJ+TJyoYz8Zo0umApfW4aT5ylZFnT4eiAYWl9U2mNSO2rzLYK8g0GN7xh6d9qyymBzURsDI2TRB94kSaANX
cwUfQGdNDpf7xB7zxU6lsks1iy6vPBLkgjJzW5M4znELilrBLxUvipfRRqjvER+vsuGgY4ulq2aX2YKDLM1hI9WVFym1IwlQHBIpl+eDxndVIefREUutdM++DyhXD0Iq
LnHKUJK6/DIjgxareYH6z84zLCah9DO4zlitHEIUDbZHxyKMXvV6rkhL3+bdBcl85yIM9OdllrMKvacu7WJvCxXrsSvDdKtKU8GJHNQ6Xy6opDvF0PAW+/Jc3ng52UPL
uNa3p0fojeKgpT7AhTDsE4v+z/HuxEsny8q6WG6duGJxXg5FDftLcyCkg7MWfkAcdGsyrBGw/nERX/VlAT+rjQQCvI7Yshk4yg9EvMXZwDtTBmoWuZy0yJa+iGXEQZ9F
hvbnU/SRD0bMd4N0IGgZ+h2ehrXbainFxtWz++B+QfwbNQDYl8jd6PssuBD75TwqC4pawS8VL4qX0Uao7xEfr7yAJlbaCENd2xijg8aRizrgC6oBDZKtKzUGwyS2ThBf
U6bgO2hzpVM70iDAxRsbW1EDGRwjfzqEqzhjMh8hEa3DThk0HSbbuy/SuJkQkbxpIGGh78VocMa2ZWDzYC1d8eciDPTnZZazCr2nLu1ibwsV67Erw3SrSlPBiRzUOl8u
8fho/Hs1HyDIVhsGVRTOMg6xtF1Am7fJ602Kwn8Q1FsarDkMbrxPKGvusIFhuDZeyijZh8LmwfiKibX/WkCyZNSO2rzLYK8g0GN7xh6d9qxJIpVN9ZhWTh3Gu6+qg9Ap
siU0pYkJE7ZGnyeN+ORRmf6UhzKBZ5Y3QfOkq5d682U9bPc/WzjtvkbrDbENBaF8YrJ/y8nMW+bp66eKMkw/ZElvTRegigbhy3a32fHRKvYvsSrKenxdB3CF8lmYUe9O
ys7XLFBiHijHIMZ5EU4fnM0lPkgHAF4YlVOrJPdcVa6S+aEI+5VK62dFyp415UjrIGM00VlWr9Tfp+3AkS0dTw1HerqyvouEU6i86VeaLyZVGWgDqyWwlKrKcOt3R3so
yPVahDH1kBucyxt63pxYJiGoB5ZjA39baL/KRjJpVzAtZhA/XJmEd9v5iU7NLblHqC8FN8TpnE/kVLIpmNKkJSTh3GDEl3tR9Ffup6lWq8hAD43LBuVfgrALprv83R5p
AqylsJLpSzYp+Qzp/Xm4V8+UsJPVIQXWT7go3UN994RWNhi82WE/OvQ+gdQ7O2WUfgSq34msx2yQHs4HH3mUj5/ntXmEZs8SNiAVj7UC6+YyvQ1z0lbgYH1o0CmLcgaL
00ndttirpnAn3FXM4UH+AagvBTfE6ZxP5FSyKZjSpCXcFvXPereLha0ka+fJfMF0aZ/Zp6Lsvleb4IONNA5vghbwv3MrNDdl4t4wD1KcBQqwTnDsK6rdM7iLc/bTqc0a
SBhMCJ2ybDMtLcywzSeDR9qhGwYQDe7POmWondys/5fxiDkdM+cksAPtG2zmL82Mgjaj9K61Zs/n+tKgzF1TpzuOFcXpZHfJle/QZlBqOLJIGEwInbJsMy0tzLDNJ4NH
dnNc9l1QHYjqyqkl6wV84mmf2aei7L5Xm+CDjTQOb4IW8L9zKzQ3ZeLeMA9SnAUKfrV3RSkAlb/j0qCUZngnGBC3sUcqk0X4YVBAc1stI7YdHpDMjYB7jreit28d+8X0
zuEezBLui8C4F4+xusvn7QQaxQBjmK5eLmqyvngn14KJFQFBXZAaDNS2JE21MW1cc+yvur8HM5Uydrh/91AcEIZDb0/HpPhD9LpYUH6T9dxQ+15j50kSN1dCbZ46oTyA
X3+j9Vm8atPQSX58HiNbhAJS6GAiHhQG50aetmf4ckiz5pIVrbLIVYOIRLAM0VapU5+FYI6zBENtKs/HrevMMfp5LibGrbeMToQJmEF7eknkaDRMoeUog81+PEF/MFkl
kkynGI6H7x8q+qn9hnbRJwe9EoO4V7KSDWdDUeTek9p7Um4g8gy77lB+uT3MVaHqMRVsyZsGCvYXcmhwVMKHK40MXsywLPH1jMspHK0EgHcoPr61vcRYZq7x3rRhVWSO
JL2OYMe7VB92zLYag8U4vn/vDKC8JelQoQaPEuHK9SFByOzABlm8bmzMXxOZOfDT5Gg0TKHlKIPNfjxBfzBZJZJMpxiOh+8fKvqp/YZ20SfbKwjCYF3b+pKD1BgmurjL
3gviT5Rm++4A+a/sW24Ll8/EwCKWOfwa/1mIAEN5t6U9fTWTUTnB5UORxJc6e2irYZMH2d7xfj/Ov90b17wpkWhmExIgztZA2Y3zQpttD4Mip4tmTuvt65r3ZpdTkk7G
z4/FGgxvRWJAkqCorzraUVG91TOLzI1t37eOa9HWka9Q+15j50kSN1dCbZ46oTyAzE+SdgQolorEIR5sWAo6B+n71tqJN3lh9VpwB0KVOhcEh69LZ3xa7LnBuKWU582z
Ll0KYRtMh3oXBBE7mfw/YuGJGG7t2QXYEwqBhedR8u3JBRGz12J4icjrkCSmGzCABHLFVZ/4K0JPhJbSl2lhg0gYTAidsmwzLS3MsM0ng0fCznSYpgmjbXPdD1ePdjLQ
vpjNG+K9GMZfIIUP2X0/ZwInZ/gWM09gKXX7lae/73OSolEA2vO23B5wDTdcbQ7fcuTIn8qK0N3kC0okwBSe/h15WmPfRu3emdX3rnYCwfsGcnMvUUcq+NZh4X9fLqTB
yijZh8LmwfiKibX/WkCyZAwokXyLKmuwoSV37jr2myDbzY5ujmgsfKZMBaZmQO6hWfe3jnp0vavBR+mSL9M9p3Db23+AHzS5dpzi+ung8YNsBNml4wijrYBmvT25JWeB
3SSxATmhWz9JM0hE/MI2wgwhyE7N2Ws9bbQhQhyY+nnHjTTItU+a52dxr3NhbBK5szG8gv1HySrvU64YDkHUZxEVBiA84wBjR2UeBofHa6o7mm92dV2DRxRwkU7Y84hG
NDzhhkKh97KQTUKhd8ZDJSjuKOktBsg797cFGUDA0EDAVSOCMVrhsgEf8qm30Cn3QXqdlAMXIWhyKuLPkpz2y0KXuxYTLlh/qoWjylghDKqS3+8BiQKUmCZTzqn9mUdK
+o7blBgkBRRRTTnID5XyUG+D0MzaH2dSOIl2Q1P5Z6zHG+H9VOaQUfwBlSJpItd78GNgkyrWLUMwvcMBAmoNZseNNMi1T5rnZ3Gvc2FsErn6xBFdtTQrAFvbiU9yRcPm
Lbqrj/1tduI0JTBC+RqS8BJrOa3n9TvCn36QSmI2cm+lCJpPbzmiftAws9x3/XX6VOtZWX881NCHQLyHUmoLg0/Txe0kp2RrQrtoPA1gcQFEb+G4V0LA/zn4kbsYEZKY
KO4o6S0GyDv3twUZQMDQQIGcIA5Fzn23HdLMoEd8h2qslUymHmIP2oMC6aOFQbjZqr8pO8feQCAZFJLhuF8wqfiZSv+dUOEIcFlKJdPmA1d9egkvka1Txjhm9vYbESGn
1icIvWPFOvLbNuLX9oo3epqR7Ytq973s7ujPc7lJ5qerLY+EoB70sZhM2SQ0CJ63gxiZF/t8eEZlDQPfsIl5jQlvrrsNY5PKmADrpFflFFmlmWC/XUjmrTqKK1wRu7z7
aZQOY/CVD59w+v2ljsRoNg3woRzySzCADOkKTdTpFoDW8+t2UerI0T5Hd7fHJkc0NpjTZ6Ws/tchvHJ4ShhZFC/Q+h6TfuVQxT/aHfMqjjxyeFWvWcP0Aajh8DmyJ+jW
8hzkm/cA9HRL66O/qFHDTsb7B0UgQhZ+IReeWjQX09fCRyS4r91md556dIENtqsZ0MB0hwYKsnGEpqtt0AingdBfgmXbovMnnFE7mlJtuJkEq05BtOyh6/vmv8kwKda5
EmTgXAbFeEt2b4OVY53dTpPuivGSePzyqMhTEgl2TiQqrgdl3csptFJbkH9n9BpoEmTgXAbFeEt2b4OVY53dTpqrdzyFhb6EePl3UzcdcKxi4vcBj0YG++JtKHtoi+CF
b4PQzNofZ1I4iXZDU/lnrDUBnEBcdeyz38v+/8rtiYW1K+anBYgFeeVItTAYv6BfNjs1j1W0KnL4BhjoV6t8mBJk4FwGxXhLdm+DlWOd3U4oKHP4WuDEpVjNn65ONQs1
PqRoa6THsk1urUBexkPd3/BjYJMq1i1DML3DAQJqDWbL8+k7ItaYXpDgPBzZNm/NLHjw0Zk/+gmCX1F3qenJHI9KVUlpVDG7VsUjiV5WJHBIsO6JCnMpzMl9PYkZskMJ
+e7PK+cRFCrP98CZvANUNNAKNE3ttfGNvXheQw5llhz6xBFdtTQrAFvbiU9yRcPmHe9aJRFJ1XL8vYoUGHMjWmJfBKqk058fiWPwO4bGZBCZ8qQbQOvM26gGWXcmmfbb
d8bRffKRk/ehjwVfW9rDrz1bi7u0btoD677HFYQOfZQ2z5VhGPS8mObytwTiiAUHreHcpwTLmPKzZAH5dgdYTl+89f+rMrqPZUTXat13hkAUKelK26qCCmqyCzuuEVgl
1OJ+v9m/2jSFwL7eFcYrRIbuNlg0hEMDMGQk2NA5xA5RINtXsnWFNN1a02OleT+mU6Me7iisvZ3IezuJClkkw5ZCItesSiXXPXCcGfNit2bSnEc+Pba0aKAAHIFrJR8K
Uu7B73QIikzIEvN1L9W/qNwo8FNwLgmRcBOo7MPJKgKoxZl264ujB7TBmJ/Nsj86SyIu35ryxKO0m7jdzKb0LlPOyxMOaLh48ZgSfBQx027Mel2t4OF5ihov5KPXrzdi
m7OUpyqr9qjffPe27Ox6As2XsjVRTqL6K+B1e2fNc2F5r0rBCIRFYWsIzFD9nI5U3sMfEMXW0idbzwZdCYTzNJ0bvupPSkv/bkE9dD0OoHKKF1q0jfjIVrNfJHZ25TJZ
8zzbe4/D5+nJBC2hE03KKM04xex6tb411BZBoYnqJLRl3banP3n94SSNDJaVwegpKjFpxnd0sN58GLwSnH+MbNibq+hu5ofyLD8URcwhm7JibuDieN6/6YLGJ2h3d8yS
FmkfuAXyiAR9/Wi1JoN0jOzIXhworPhL9VDYLhDefoBoyCKRb1mFWWnG6cfL8fHHmXwj/171m30+XXC2NXYdVvVSZHX5HTdsJmh5oGBGNv9zvtNdWKRitceobBXNnTFY
AcTvF8gwooMKmKArv5m08ILWWp/mb9HUcy+dpaDoE9Q12fsN2rY0eJ3Wps9zpfATY9Dcw2LKdkS3YveFiKVikR5Qc5efOrc0HlGoJdu1n0Zl5X2RBiZte9dXW9FxpC1V
bEpWVUfh4NbUCHVH+8Jg7qrH5aA0KbB3VBfMWnlkzzyMoz5RX/8njkCDwpxoq7BtCc7EdKOew+mX7J/NJc2zEKQtlgvq5Hp/YwOX8NE5+nmOfyoitHTO23+3q4HrZ2re
TcFSaIX+D3Vr9IKYPjM1YvCaEpwB1mlMLklc5+Rj+iSwY2CAOTPBB3Ej5Ur7qhKQdYc3Q6PCSJCGMXuYhabpaRY8++eKGT0NNhrFlV13z9ez6s4HvoNtgafnSWkCbwbA
CseZ302fZ4vGrvx+W75VR5H14yl5+T7YgCeilbofl+nuBRTWf9hm9kUvEQr0tVrhRveogmJ/63sY5vjruB6VsHWHN0OjwkiQhjF7mIWm6WmRZm8hXQmA+VZd2DcRb8Dx
961Kjjok0iHYUyDIOR1YrmK0GwRhCLDGcoq8CONojggJIum1eOIKoxSiV6VuUAFsNfup4EtVD5o50Dg1MI6e/lOjHu4orL2dyHs7iQpZJMN32Zf+u7IlcBtzdOyO338N
0pxHPj22tGigAByBayUfClLuwe90CIpMyBLzdS/Vv6jcKPBTcC4JkXATqOzDySoCIkgqXbIddGPWlhDlt8asgUsiLt+a8sSjtJu43cym9C5TzssTDmi4ePGYEnwUMdNu
i+b/KD9QLEHxTnVA9jBidZuzlKcqq/ao33z3tuzsegLNl7I1UU6i+ivgdXtnzXNhea9KwQiERWFrCMxQ/ZyOVIgH15Dy0t5sXQ8q/6/jy+ydG77qT0pL/25BPXQ9DqBy
ihdatI34yFazXyR2duUyWV+TM7Q+GTBL2TjgV9wllEHNOMXserW+NdQWQaGJ6iS0Zd22pz95/eEkjQyWlcHoKaTgoUhKFQBCMV0T47NkJjUnIhGlVmCEUtem9aG98kDM
Ym7g4njev+mCxidod3fMkhZpH7gF8ogEff1otSaDdIyuTmZkAR+X7AxFlOhIjI1waMgikW9ZhVlpxunHy/Hxx5l8I/9e9Zt9Pl1wtjV2HVYw0f9r9iO5xyWBPDEbzGlJ
c77TXVikYrXHqGwVzZ0xWAHE7xfIMKKDCpigK7+ZtPCC1lqf5m/R1HMvnaWg6BPU9DGAF5rlCG6vax4DTlblEWPQ3MNiynZEt2L3hYilYpEeUHOXnzq3NB5RqCXbtZ9G
hHsxA6a9oFJCPaBN9AjG0mxKVlVH4eDW1Ah1R/vCYO6qx+WgNCmwd1QXzFp5ZM88OPg+9fzFBdKUmbsrOqP7Ldh28aKDEf4rLVjBA3mz2ECkLZYL6uR6f2MDl/DROfp5
1b/jVxkm1XcE0wSLexS16N7ISDBUwEduHZuV1TtCLIzwmhKcAdZpTC5JXOfkY/ok48tMwLZuIDE2TSZaZWh4e7WAk3mtmQzRuMA4kuAotOT/EpVm2t5pDH+0KaXMLopd
o7htMM8El3e9MUu5iBP1C4IiIzj12Gizte/EMiWkchLkoEDaV9xFGpQmP31NLv7LOWQXKT7Tbs8iCPlhnTl64X9V5lnijLjFn4O8rkIRQ2SkLZYL6uR6f2MDl/DROfp5
jn8qIrR0ztt/t6uB62dq3u73aNIZ77ObUr6g136N6gjwmhKcAdZpTC5JXOfkY/okcD1fqi8OcQy1US/UzandQnBu9ZZdFNZIMbh6monbUE51BIt6OZ2/Nc3aBxtP+J49
ldRpmFpJMe+zMEtg2kAf9/hAOk6p/EB2X5niKfp+s46FziNLDMOyrZbx++vwUaAqMbZ7uFk12HCJ6bG/2vpDfyjhkCKrExg8IgL24ttT4SP9CHiOj9jb16Ag5NokpBFt
gF6y6gR2QR8DRhimIFlgDJVf3v1U6mtnUXtso0twlZDzqW/X9KkQlHFPPWxdWcObi6qCfPbl59E4T9U0ypw7G3u7+YddZzTMjG6CBHCb0D4oyEHWZ66gIV19prT/uaCQ
OuyoWJMHtqc9MtgcGSly3SFNCvIk1vcwWwnl5a/LEwIpPxkKLSoPQSOoXO8/hFKsSAqCKHHzEitgzg+VZX8Ji32OYm3Jhfo+HIeWKtqcIYf11GMdGopG5DcUCPndfwUw
PSmVpocxbd51mQts0+nvLTvtDHXdZZPhr/y9MewweBhEd3RY3uynNGRCkFhc3VVMV3NIB+alHGbCZ1oy1ix8SmyW1DlA0ObAbscTvBZ0p4I2EgoDqnCEVq20+kTLAwXk
65b1zQLKVxzCyixDX2+xEag55HzDfftJiOilsTVEMcKrPAGK1Z+zOb0GHo9vvU7KD1WLPj8VWPN/YRQrn7VvTJm+Bmctkk5caele0eGG1xd7xqCUNVolHb1aY0m/p4+L
jwZTsdSxdVlEgGlr52stpvXYwCP5ycrAE29XFqNE+OM67KhYkwe2pz0y2BwZKXLdJGQBtRhAu5LbqsUBhdusUuIUt92boHRyqYz7gWW90wr1zjH4IYPBIsz/+HYC7tZG
RPMe+Pv279XMBQIE+YWNnUd87EmNEL2/3G52zk0ArWDiFLfdm6B0cqmM+4FlvdMKQnVO8QGklFUvx0gPj7uvYllp2qygc+ceAAt5PtJ/uZ0273KEDu6reo2UxFqrNDLv
xnNbuW5kP1RKCGGyDKRH7hMgdFAaDjwCoIv/YIBSP4xE8x74+/bv1cwFAgT5hY2dEPLqH+vf3s2tDPsiRv1lWQb3ZNu0dahRkx2LmDqfb9IMHDjclz4ZJGNPRl7f5z7v
Cz3B2Dzdj9V1C86J1IsPlVm8DR2AzgdnptgR0VimOV7N5IGhVpJLZdtm+HbhjvxOD/H+1EI4/wBP/PTSFnJKT+WArLg2q9ghEGMbvLugViaEO1LPhxGufbY1nrn+AM2x
GpxsbRivgYDw9BBeLrwJrJAINtUfIQnmIvrH1H6Sk0txoBIDECt7ah5rfIQ9HiF7zuY+X07c17gsgSKAmso3J8hTLelX4usEUHPkCWmbw3okSPfYy8NR2c45zDNXvl2s
EbRqUdVkxjnLixPksXPk/klehOCcgFc27IX0Aohmpyg/9/urhlfcwmT8NZ/CbZMKzv5ocQ5w78VGfgs2/okcI8jp3U1ukNsEILyE8Ndfb6yJOC4DhzD1tIrZzjzaaXzT
El0ZcBS3sBjoznWGhDpCLdWy26WATr95Yxz48zi7vsbe4/cuRPcoQ8/e4t4rIKbAO+YNFqCbauHAUqnyP2q2/84GPm/EctVAbBFDBeyoJnSohOM6oo3abLT1nqEpgKaI
wPI3y+jVzDQLgAHdlQEPFeBaydVJWWabnj1pQb3XuQq13XDF+syrjmz9q0VNHiZZpBOqLOnMBlNjVe7ary+SZDENTq2h7+zMrm4UVKp5ojU3+rGMupYp13FMtvXTZ+0h
xymw+FMgzQTO0olNl/pvCr/2P4senIOwHeZhSfqfReSxpD/5MgxD3Lu0e37P72VRpo4oGf2CaKyVKzSlGKQFbH50+v6IElAJ7IwO3GoGvz15ssf2iKXJzedtWdYsRslt
xEep0dI1Myezwdyas1d+hYHXt6qX6M1ubh1yezaHBcwBOiaLivRq0H20uIOJWbehoqY6uyyaRB0MwtS/iTEuSgfJUWQaHgbFmYkzumy43DJgsG4e6ywWR5VOJsXYrMY+
6+PqlF9kFRc0e9hRZ3/LciFcsI6OpCyLM00yxwi8GIjmYZrzgb/FN7VovGbra5Y8wbdYdBjuBf/5uACVYcMApPBqach14HQwjaHBk/Hmu/qFs9lWHIn9XckN0yAEc0S/
XFJeDSOMkUefAAdciLTlSeYeHx1D4H4W4eogllbcqT0WlfrkUrgIOowvWjGBjWrxT+pYENSLQukftZdMz0REAEHQQdD1O/BFa+56rVchl+14UVgQc65mLsvpr+7e88bN
z1BIR6+qMgDEYjP6eW5e5GcWPM93BzVP44jjI4xjzZSVzl23Ctzp1tPQ8b4iDv4X5mGa84G/xTe1aLxm62uWPKDmpa/6BotDfDM66i0xmzCG+s5mfc0Okp0hWcZL1pkJ
GkO/PUacvdGwVK6um/SvRzqYcAEy7WgOQtBKCKCtVfTEu49H2jd6Boc98RxCT18aUPteY+dJEjdXQm2eOqE8gGRcNwQ7ub5FuxILF2M1GMo+PYucVyqTCRO1eT6FLOcK
yFIJ0vGGnoJIZqjLpNsHTvqZZlFlYw4genZZ0Nlt2T1Jb00XoIoG4ct2t9nx0Sr2pCAt9pVb3CKnmXmRKqwKCVyjLI/SgGYlGNtDvJgATTBvKbOeAsxbqKCOf4IzOd5z
U6bgO2hzpVM70iDAxRsbWz2UHhRP5OuAUuUz9JhC5sA2YCEAUJAJ4riSwfLUO7S5KUgh18wfkkV4Tg5Z0+FRdV2BQ3hgz+JUqs23J4GHjwqwSoavkXA3OHZVG/s4ebCb
6tP7xeAnRkzZM78zvIYFD5oGCa5kSQBKDk7N9B5yBeZX/Yr4Ly7ww+MbVhLn8Pt5SFoFHdhbuBJKUDu/RZf25b4dXkPNoMohK+g4PVmme82olsw9OOEGMcPalLAav+l0
MZ+AW6CuIynWQ9SXnhj7FWTH8Eok44ZMFr9JoAfhyQlOPVG3GcGu4LQYz/Z/Jqj5RbM4khcEkCCDDzYdXg+Ww2Y8PWKgmmFxlZ76SCggnGhYojP1D2/DHhHjjZNzdsmv
vfZvvPJSmeD4yVS2niuR2dchdOHU/fp+Zqxg54D48QTglfNIJbrLB0nJlNhMVed4V/2K+C8u8MPjG1YS5/D7eWq8ZxKOiwT2pg1vzdLh2eS2t9evRLSI+bp2ZNET2bku
v+TnZzKxiZGKq6R0TUkR/6QU1zt/RUHSGcep8OGwf4aNtsmI8HrKLp+Pbe/vVbZ36ODut6g1V6zcP7HyYWxacfetSo46JNIh2FMgyDkdWK6I672xoZ6KsI6yXKdB4e63
QXd87gim49GRkF/kOuLDVVhn7rca2mmehrW9BM2crGyEcr12vis6tjw5FMd8mNW0e4RnXO/bGqRwV2sweD+jFNt8hy2pwr37UeY8AMqLxYcju6iclLDVhD1csYe4iNj8
OX8WZCK2w6CQJ0zJSgKJIwwJfhToQm19bbh6ht1geBW5833Ih5lMC/sm6ONF7fDZnUoDuJtE1C1TCD92i4NlO58FmiTCF90lCl9I+aAv4YHmYZrzgb/FN7VovGbra5Y8
9n+agCTTLXVLqtrOiPvSzPah7JpG03U1RWgPwGmyQRdYZ+63Gtppnoa1vQTNnKxsjJVVj2PYVCelDduba0JxJXPY1zyWmWoz4ev90dtAsyc2UOtyVY2zRYHSzPRD/6pN
h9tbdkseeC0BGXGZ1tcUz5oy4EAYEQHbF44acxKyKPMemc22UD+XnPruCzdRGpdls+rOB76DbYGn50lpAm8GwH+FMLSjBDHvBfMNpzRWIErJHfFUxnZqhf8lD2tmOBPQ
BubpSVSy3vWxe4LrmnIlggBvguSgMmD/B5OfvDWwVmdl82Ul8xzW6v8gBiZbo6o3eXrLOFUuVxe3GKiGQHSH85TPSxQ5OV3pn3j0I3adBYgbg1M6qcLEUYvHHwmWzrYx
Rm8zRLvUyoKOl2L0/9WwCpxxg0mo9YQFRpeuQs9iANSlXVkqP4UXnQkS4x+SXGkLrgsc2Ga+1k4+nHxPzNf6HmJu4OJ43r/pgsYnaHd3zJI1izEU/mYxt8uagxMVxruq
WLEltZ/nKkvHzJEhgE1BiuEVeYBtHot7eYFbO3lBiAEaQ789Rpy90bBUrq6b9K9HOphwATLtaA5C0EoIoK1V9HcidPEe7appIokgVYjY+aeAHY5DNWTQxzk4ttkDvlZ4
lbuS/Ll3tgwGii4ZN5y4h+BaeliaO+GoZF9REHtFsswfEoAUxybwdJIP++JiF2ePy+/KBcRvy6e+qn/l5K8lCmRcNwQ7ub5FuxILF2M1GMo+PYucVyqTCRO1eT6FLOcK
zkT7gE6lE0QjZXvN/sim9USuqtFaC4ssy+ITOZpmGMeSdyHHWSST+2oZzASxm0kZ23yHLanCvftR5jwAyovFh4pF3VgqZXG128SEw1ZmpPNErqrRWguLLMviEzmaZhjH
CfIpqd6jc10/HLqSFXX8D8ukrewpxK97OhV9/mvf4zVc87IOTcgLSaToZt+lYHjUKjSSNhGh9eaWp2daon/nCaJImbzO9LDNZGsv/EMA/Lu0PRx6aK3rXdIIm1whlJ/G
rDCutQr4IPdJScvIwlUBQ/etSo46JNIh2FMgyDkdWK44xfmj4SZ3Id/joEPVC6HoQXd87gim49GRkF/kOuLDVeciDPTnZZazCr2nLu1ibwvjS3BifyzZcRp7QOKB2kcx
S2WVz4aTVE7OufJA/URcRhs1ANiXyN3o+yy4EPvlPCp/4U25pCQPg56TFSw8iK10hp0YNlt+zKnDnf6GRmoXuQHE7xfIMKKDCpigK7+ZtPDJxXq1wd+URapXjhceQYj5
f+FNuaQkD4OekxUsPIitdCPKUTOtCxhqvKbMCimya3EuFuPfOTpbIeF/OLms5p5dDlnCS4SR+JHwqj0zdMRHHWRCrLYr1iNl4IfUMQ/Yqv4YGKFUHp7gGOm6D0t0MQAU
JI2Gyd5auOfqhwueZ5Nin+vJBKP6AZtMHMHYlkijlIWuLO+vk5M9FpJrEpM5cq/x4lNnQHEmBf+QPGwtBpFO46RlDZjV81Lfsfg+OwawMp4Uj6BsHiAw5ImsfPvTOIZc
B8lRZBoeBsWZiTO6bLjcMs0VXA/QfsMuB7uceA/b6GhR1K6352JQ5BqnOT0FE6XD1YpLq2mpR8mah8Ho/AjPHKK7FTu+CiMspzG8gEmtnErU8IuaO2coOXYq1/cKXJDf
v5VfjRk5GHeULvOYmkH0dDOOX/co2N40wTFr6Ok3V734t3d2NWFmPKU54mamTgkJX6WTdttuQyYlims0HGLJIqoVzhcfMaHM8TLruaat57+Fa6f7/DwE14gCBA1xXKj4
A/Oez28fJyZqKeaz2FZdlTaxS6D+sqZEClmQSFVmZs74fIioM67EveIT9bMvhFXNXUKMcDSxK64sxU/pej6rf8cp9SX21C5UIiDEUSF9x3q66zcPOYUYIXxGEnEkKHQD
+cfp1QatrPshrgZ6c7S2qG2jnq3DMPzQOUM4z/T7G6ICH83vxX/QWNq//2crN0intKTwGhGAMnThi/rRMbVyvcW8nGuEK02yIiYQwuAhfp1DHgvgJucXol5d2YFlnrsP
BQ4dgDIp6l9J394i4frs7Ph8iKgzrsS94hP1sy+EVc258ou3qJh+2NSKXI86f1Fo6nuZShhJHfH60fBGQcSuLzxQnJVoIcyRPkZ279O/BHgrXdGiKqO36d9UefHi6fsU
NVHAyhDll5eFLNljKEoqf9nBtOOx42LakJrm6DbKcmUh0aetyYTDNp9CW5DPVtU4z3UnmUUaT+av8JazJxwqaqdfV7w0VqyWxxkIjqblWd2i2kRDfDS2agjeG8kd/Otp
/lFAoxmldu6uVRym9eqgIn0DgrVm7rXl19tks2xBGucgCit9mBHTsrqGvLMDAbRZ6dxqNIHlH0MGjeqpG0BjKWutIJ2b2MkefXUP/lAXoYGiX1vgGnK+6RkNEDk7n1cr
2ktNgYVQxe9jrPB280O9PA8g3pQzG5XCf14bcQDjt/fLSpeVVQNMW3ZBW7zjh6bkpNF6HciCx1nYyQoUw+kKfIplx8KUWpOknMBrGaeLhLsWmTDHZnCMd7pnCvC9IPQ2
Dp0gdAh+AU3pEgmPgE+3iuqpa5ozQeJ4O6FKxGTUHEpnxdgNYKcurSLoAg4DdLLCiXUQ4+Cjc9bUEic48mT7aYj+41bml+OhWPwdisz+wZplTYMmUY75B0TTk+mJYs6q
hAFDd3gSD52jt1NGm+TQPrdUlI1wZaR5Cbc7PjvqbIES34Nv7MUUhdQ4C5bZaH4mx5EzGi0GUCUeLzCytf/454bo0DIH8eQPW7hojuewM2kEZGrQSrEwO8JTEm9xBXkT
u7CqpPScOO98bOm3OsXPizomWlv/r0hy0mBV2cZsmWzDqPHGSsNJzA0QOjAvIv5rRadI6aAQke0Uy6V1oQrn/Vze6gcPXpZdbwVQdUrH9T5tE9yyevGUuy01rHBya6rX
4rff6aK2gF1OqpTbmaxyyBGXdooJ1mMYQB8ApdwwOCqL0360y0qrLdF3Bb9iRzne964mA0tlkkOnmGtUkQVGTOizszmZ4J/lSYwY5tnM5LDBDYR8LHGHIIpHRkt7FGKJ
YbPV1Oa6tMG5dh6MRu8Rn3ZvGkd+NNJUctF/cjpxLGg//aBI8k0MCXOsz5twfu8wEDRcuZcz3ZBASUEugbhAaV6ye5RhH/VmJK618muB3ZsSEYrzKpw7rhnux2WmtWqS
x8XH7NEp+xPv04NHxJhWfWGz1dTmurTBuXYejEbvEZ92bxpHfjTSVHLRf3I6cSxoVfDJsDrir4TnyApuH18pH7uwqqT0nDjvfGzptzrFz4s6Jlpb/69IctJgVdnGbJls
K2XxXHeoibXpdihEW+nfCPTLtuE9L0HrqkwxIWzXr20LyrShRnvTy5qa6oR71dvXxGkkPcc41D0feq1dZi6zuLnZ2n81hIaaK6XFIp51cAxmADq3HxTURtS4My6IfO8e
IKoLqRA4kPlyd16kM0A6VhSNltGzfHwrJjcsV7x3S6wkmc66dKLIyLw/OxjgtWXzKAlN7eKHCm9zvqakTBrIKgOo6QMjK/tEfF/H/nOuznpFkLcdhCIw0bzm6JONWLkD
JJ4aQXGEATMuL05UOVzqrdSsfPeyhymDSNuEN/EBX8pygqWMCH7an7xYi6SbUKjF829ez1zl/6SfIOLaOfUCiKV6rUiLohzYG7duCZ4BIEAU9egoVTmB0tPpETx/nGmP
gvUfbULzbxBVb5k22nsmZXEzODspEi3lTS9FPLXjE1JU6hWESvStgAlyL4wp+WeFcoKljAh+2p+8WIukm1CoxfNvXs9c5f+knyDi2jn1AojrPr9zRgQcvEeCxybF3No3
C8q0oUZ708uamuqEe9Xb18RpJD3HONQ9H3qtXWYus7g9Bk4qvWRRp/4GPTyQWGH6O0PeFS0bouZ5usIIK7vyiHZvGkd+NNJUctF/cjpxLGjaG2GOkHDb8SGsoBODOWaY
yoDb7QwiqZuYOqt1h4Bx316ye5RhH/VmJK618muB3ZtKOnv0en889Wg7ql/GxkNuA6jpAyMr+0R8X8f+c67OeqN09YI0rlsEsQ8t0sc12EfHTFJw+LPEr4hvv21cW3aH
zPe0rVq2Y8wJ+KauqKmpSYYDbA1/ONrOsiuSL1VkjHgzH/ygnPDqG+V2iqch1F5b2Z+Ozm1kSdg57AuwcvHmN7uwqqT0nDjvfGzptzrFz4u/J0rrrGC+n3ZsswIUur+U
kOTsAzMety9X8U5yOmTLQUWnSOmgEJHtFMuldaEK5/1W/I5zCN1nn54rHTN0MQ/YFgsFTocqq5/SF4kliYu8+rZyDo/7QDPwsNKGCv9Fyq27sKqk9Jw473xs6bc6xc+L
vydK66xgvp92bLMCFLq/lHVtuMfsg5iBBsnfaMRQM7F2bxpHfjTSVHLRf3I6cSxoJmF8MNkcVCvylJLxz8lWJH6bn610NsI6gxBhsWDk1najG7BkF39ky4Idk/MqFgFN
829ez1zl/6SfIOLaOfUCiHzF/nCkIT5EYZj5V83CTOwU9egoVTmB0tPpETx/nGmPXRZ5E1KPYW29PRm1/BMUWxO2xPhrkVujBCST98FAF9HM97StWrZjzAn4pq6oqalJ
0sYUzH0WfHcgZggLefeKdbnhVJD4zGnNLPy7dqIRpizit9/poraAXU6qlNuZrHLI2+1g+sRAyOdFKhiqMn1hHr/QNhiwBT7OTCUgCittvXFMFVZBLu/YUKgr3fuS917A
C8q0oUZ708uamuqEe9Xb1zizEX5uaLbVkxBx6CpRvKun73yggvRJNcK3MocvkHKiZgA6tx8U1EbUuDMuiHzvHsCQBIjok16yIqFG77G5l0OFAh7IvmrnFctQeOdjZ0EI
TBVWQS7v2FCoK937kvdewAvKtKFGe9PLmprqhHvV29f9qs7/hFX7/ISIf8KlOB1vRs/yfOHCGO78KdV4EmEc7PNvXs9c5f+knyDi2jn1AojfUO6EfPIqlGOZtL5QhpXx
d6lnp1xe+sHrMUBQn4fRZLuwqqT0nDjvfGzptzrFz4sKSlB6XcUWjp6+dHwxsnVUw6jxxkrDScwNEDowLyL+a0WnSOmgEJHtFMuldaEK5/0nWzk5hhNAyUmAClN3iJj/
bRPcsnrxlLstNaxwcmuq1+K33+mitoBdTqqU25mscshJdeq9XDNapaOWlIzNvxjci9N+tMtKqy3RdwW/Ykc53ujiemt+tiuj/okSYslm96Xos7M5meCf5UmMGObZzOSw
BU6M3VFDivCStkwOa6Ey6uH8c+0z3vC+0sG7Tqas0yx2bxpHfjTSVHLRf3I6cSxou44U6lP0n7YI4Dg3k2S5uBA0XLmXM92QQElBLoG4QGlesnuUYR/1ZiSutfJrgd2b
CT1w7gPLkZzqmX7fmJnnepDfoxc7kZvqrvpSSfdYQADh/HPtM97wvtLBu06mrNMsdm8aR3400lRy0X9yOnEsaI6Y4E1rV09ii0ojjzNIJW+7sKqk9Jw473xs6bc6xc+L
CkpQel3FFo6evnR8MbJ1VCtl8Vx3qIm16XYoRFvp3wiSFAS9yCzw4P27JtD+FJOdC8q0oUZ708uamuqEe9Xb132rywOFoOidSL3Ntxj5sin7ONILQlHw+K60tJ57dfo9
dm8aR3400lRy0X9yOnEsaDpQSNrGuUSTVjao5FRP8GwrfmIU9Jdzpv2kNypQa7dFXrJ7lGEf9WYkrrXya4Hdm06nvi9x1Vrfr5GHpc/AqSK7sKqk9Jw473xs6bc6xc+L
rtE2fXoXrJT+V6gkVdKcE+izszmZ4J/lSYwY5tnM5LB9mQQaNF2VqgIjbO4tPmSNIohYYKcgCV8X+hB13tIyn3ZvGkd+NNJUctF/cjpxLGhEGT2vlfHy1d303svB3uWR
R2QdPZmMoCnZvfQY5mC0SvNvXs9c5f+knyDi2jn1AogfNl7aDHfT7rtjh6Ke/EKZGpJtX1q4df5Oeu+VaK7L6biZQPyhVYsSQcnAQlZzmAJqxp7RKs8+ohSU18s0XEzA
rFkcjcMWOkihYDoO40u8DBA0XLmXM92QQElBLoG4QGlesnuUYR/1ZiSutfJrgd2bZJI9XXmhZ/EDkldxeILElNZ2PS8H36DETzePr5Q/YLkFoQKVvhZ9krM4qR8IyaGu
eTLNMbIKKCScOjn4/1Gge+3I3DKhEz7Atndj2Yj9C+YHxbbeowZma/w4VaymQicdZ3JCNYv2zsw6O4Y3Fh11pzmSDmgE1eVmmdPvwFH0mvqeZeG34SZJpchBm0gBeLBO
LzJqvbbAIa5WWAWE2ThUrbac7MX0YFQB9C70AlP0sddo/XMu18WpaxOLy37JDrN6QLfcNwWVyqlTPFJKx6pcOfWcpMOkZ9FMsqlVshjR35bO4R7MEu6LwLgXj7G6y+ft
1kDeTQSet2EUifMY1sn83J+onRTU43MhnRaHMYxZTbJmaL5shwKiUv3ag3eIrkjLMgHFqkh94UzSzJFAKmO3eC8yar22wCGuVlgFhNk4VK22nOzF9GBUAfQu9AJT9LHX
WM8YBGWA+D/f+MlxVQQbTnKfQQHtbWd6JzZFTulSkls8mJKn9NqaY6a+XdiaqLG50gaKrE12QXykuAqljZv9e8Cd3b84K5sCXKusIxcsYqo6mHABMu1oDkLQSgigrVX0
xLuPR9o3egaHPfEcQk9fGlD7XmPnSRI3V0JtnjqhPICHWZVFN1C4ZdsqpdxEhvEcujfnf8LQmPdlSAnpAsgap7qo4MVa0I9vRufFLah8e6yZ5IsQlnZu5HCRPpCWbGfy
UPteY+dJEjdXQm2eOqE8gBwm8CG/bTCu986GrQQLdIVcoyyP0oBmJRjbQ7yYAE0wbymzngLMW6igjn+CMznec00IKbotZEpA9PUzJR96LYN72XigU3os0LOR/8JhPjqQ
KY1Zf/fpHuB+t3HLe8UeLFnmO+PbE3TAGISJkI4tzZVhUqSvC6EjN+JM1BloexxEbNjANMVb7cV9YcDBKDW+lawwrrUK+CD3SUnLyMJVAUNrMv9rrkdKLz2mtglJWtfU
Qd2Bsr7M/XrTHqRJtKLLdTd9+ykY83thG6CTCcgYo597aNzBUm585CuDtg+hffA6YvDwQ41FOIIpXBM/WVkmlcWLmIJFAjV9f1zyAzuGJEaRhYrmuGDgXzhGnrKLCFZb
9ukvOzjIEB9CuRM8DHjG6/qZZlFlYw4genZZ0Nlt2T1Jb00XoIoG4ct2t9nx0Sr2vJdcdnOwFvi4cs4HGTkYZWTH8Eok44ZMFr9JoAfhyQl4vqB2mLnyPnW/4U6WjGOR
DlnCS4SR+JHwqj0zdMRHHW0dJMul6zgeHMxKJ7hLkYr7DdNTBouIDyd+0h5pIKvK4WOH6gw0EEVWFWmXN83GIcoo2YfC5sH4iom1/1pAsmR/4aaKhKCs2VK5o9wAbS0w
5KlVqk9tOd5FRo0v0sUV7LOtjYKeg6I3dA6oAZkeB9qG+s5mfc0Okp0hWcZL1pkJSzWLLq88EuSCMnNbkzjOcQuKWsEvFS+Kl9FGqO8RH69l82Ul8xzW6v8gBiZbo6o3
eXrLOFUuVxe3GKiGQHSH8yo0kjYRofXmlqdnWqJ/5wk+t3Gadz6l4NKBsDP4mNCkOphwATLtaA5C0EoIoK1V9MS7j0faN3oGhz3xHEJPXxpQ+15j50kSN1dCbZ46oTyA
i/7P8e7ESyfLyrpYbp24Yug/F7xFB9nzv6lCCwg6vAgk17i51Woyz8BSdOirele7PJiSp/TammOmvl3YmqixueciDPTnZZazCr2nLu1ibwu9+xeoVq+1A0AgS4AolYmE
gMjrZpglksZBGY2K2V0OkJUoVoCc0FG5zuY9it+Z9pg7yEf8Obx9sNllv8SVXJcLgEuAcW4dhWYY+VmVdm0STSTXuLnVajLPwFJ06Kt6V7s8mJKn9NqaY6a+XdiaqLG5
VdmgwS2YE7P6+awFzsnab6u3dUBInu0gQUvkuP2C6FFRis/HcgmMcYqEcrzgLZraUPteY+dJEjdXQm2eOqE8gMxPknYEKJaKxCEebFgKOgcpjVl/9+ke4H63cct7xR4s
WeY749sTdMAYhImQji3NlUwANvdA1T7qnx4UPedeba9QO6P0Ffi5bhAiJhKTLw++e2jcwVJufOQrg7YPoX3wOkbxtkYKqN5x7+D8WK+9SZ3CIvhpwr2w3aHn/lnuISlq
dKDCikEGhwhkheGEEox1RQajbUkpjAwSYsCmNPzWjApiXeVoE1UCtMvyV2b/jx1lPTCOW0L6tA0RU/Uqf982LmmN0nnB89mfsgKZ6iLhBPjuXCgsT19diSEZ0EZKsN6S
BubpSVSy3vWxe4LrmnIlggcz/AzImCCIvXvC41biajt1wLoUYjnAAEjwaCBgCZ6KAQVYFhZzpR7XPEeXoFshVfWcpMOkZ9FMsqlVshjR35akLZYL6uR6f2MDl/DROfp5
bvCeJE/H4vm/Prdm0oN2W1zzsg5NyAtJpOhm36VgeNTi/GXD1i4qS8XAKd+CVfX2DmlC5SuGORuXNB46ezok/p4xufjI6B0gc2mygOeqA0devPCGdv8g8eLq8q0NYH8k
1kDeTQSet2EUifMY1sn83B2IiiOtclMS7WChCy0HJphHg7h+EAMrj85zck+SKps8WZreS95Y2M2X/Wl2rqStzrac7MX0YFQB9C70AlP0sddo/XMu18WpaxOLy37JDrN6
aIAT+6h2/ykPNL9POFEc6vwK8Uv2deupdm8CKghvT/urpY9OqzrTG3VR9UcCk3LYnreOuqgKTuhm8gA8sOhYIWrIrzzIZ4liGaGdfJH4hNFyn0EB7W1neic2RU7pUpJb
q6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCGvq9BUE9ehzbfKMJo3fxlAR4O4fhADK4/Oc3JPkiqbPFma3kveWNjNl/1pdq6krc62nOzF9GBUAfQu9AJT9LHX
aP1zLtfFqWsTi8t+yQ6zekC33DcFlcqpUzxSSseqXDlRxaX12eJ8e66Eny/lQa8j67CtcLqZhKaAsp8/23T0oNZA3k0EnrdhFInzGNbJ/NyfqJ0U1ONzIZ0WhzGMWU2y
Zmi+bIcColL92oN3iK5IyzXRZklXN90yiYtIgfyam9z/quZ2O1gb9ksqyxwSuwFISNZodRTQofIbQ4VJyf6YGbLhoGOLpatml9mCgyzNYSO/gSrnhEeKVPxiHcah7sjI
lM9LFDk5XemfePQjdp0FiFDIArDnXd0xyUa9txiQK2d6XljQW/w7Z13IrwbcKGlnyR3xVMZ2aoX/JQ9rZjgT0Abm6UlUst71sXuC65pyJYIHM/wMyJggiL17wuNW4mo7
dcC6FGI5wABI8GggYAmeiuCzNy12oN6Efmw/9Zr49v08w6jq3wOTZMa4vsKf8Aeys+rOB76DbYGn50lpAm8GwJF6K6HHO6xEGgYSCov2nhr8CvFL9nXrqXZvAioIb0/7
q6WPTqs60xt1UfVHApNy2J63jrqoCk7oZvIAPLDoWCGg5qWv+gaLQ3wzOuotMZswDgKDvunBkPGBD5YQrrZlq/3DkbC/vp3zYTAKcp47CuMskRGp4r6EAsD+85IESFm2
Ym7g4njev+mCxidod3fMkgHev26XTDn6WRlCS/zCYkr9w5Gwv76d82EwCnKeOwrj+0Apt/o1NmmnpdUMmlsP5Ko0pdXPb+FPS5QPQ0nkscfKKNmHwubB+IqJtf9aQLJk
NGLr9Dv6aNsKKpa1QaY2rP7hwC69Jj9XnwEMTFkYw2w3ffspGPN7YRugkwnIGKOfrAvuv6hQ9L8wKEeFuogYxGdyQjWL9s7MOjuGNxYddafZg8Goa19bmST21RD1oNRU
23yHLanCvftR5jwAyovFh4pF3VgqZXG128SEw1ZmpPM9MI5bQvq0DRFT9Sp/3zYuJ78AR7LAQOx3rnlvExQ/brLhoGOLpatml9mCgyzNYSMC3PSzoHsREGVPfCyYvLDk
0eUoUSJfeFLwbAtTORSZybac7MX0YFQB9C70AlP0sddYzxgEZYD4P9/4yXFVBBtOZmi+bIcColL92oN3iK5IyzXRZklXN90yiYtIgfyam9z/quZ2O1gb9ksqyxwSuwFI
W7z9J3VFbg6BYeC4mcQjykC33DcFlcqpUzxSSseqXDnbfIctqcK9+1HmPADKi8WHikXdWCplcbXbxITDVmak82FSpK8LoSM34kzUGWh7HETKzWbxK0/Nr737CdKxe9oP
5YulsJuxllqZGn0v6sEgA2sy/2uuR0ovPaa2CUla19TQdl1tmMAI7Sm/8no2SrttnmXht+EmSaXIQZtIAXiwTsy13KeJwLIbOoWXS6NmoT0sOMGJXF5BSrRjaf1nmXIw
3oDnyxaoQmYjvd/O6p0uhHMzpwud+P24L8GtEcqTGb20t20pfGoquWW+SPmiN9yLdyJ08R7tqmkiiSBViNj5p/rscHMSSZCejGsP4cxCmQHbfIctqcK9+1HmPADKi8WH
ikXdWCplcbXbxITDVmak82FSpK8LoSM34kzUGWh7HETKzWbxK0/Nr737CdKxe9oP5YulsJuxllqZGn0v6sEgA2sy/2uuR0ovPaa2CUla19TQdl1tmMAI7Sm/8no2Srtt
N337KRjze2EboJMJyBijn+xhGUUlL8YR4IClV7/Od4ucS0zKiohbbdnA46KuXpTklzc0FKeNcAZw4/6s2Yq8YFMArvqfdj1OM1u4OuwLpvq7gwxnEAqsMfR4KW5bE5X6
9s8oW7v03dmaaynex41gDqo0pdXPb+FPS5QPQ0nkscfKKNmHwubB+IqJtf9aQLJk/vGWjfFLXZkkXEggzHcsbXKfQQHtbWd6JzZFTulSklvkdXE162C5zftMeqEG+T4g
xUndi6LOcsGgBn8zknXvH4fiPagCx1A1I8xpQ1VfKPCLAiJzN2BVrO3CiUB+cH3jruwWJlt8+GBnPhaJFH7eu85E+4BOpRNEI2V7zf7IpvVhUqSvC6EjN+JM1BloexxE
tOedXE4YVHbUBVL6kf+6o1MArvqfdj1OM1u4OuwLpvq7gwxnEAqsMfR4KW5bE5X69s8oW7v03dmaaynex41gDqo0pdXPb+FPS5QPQ0nkscfKKNmHwubB+IqJtf9aQLJk
/vGWjfFLXZkkXEggzHcsbUqL6eb9UPyHPHho0lUh8eRevPCGdv8g8eLq8q0NYH8kJSOqmHfq4/01r8uJCDDAR3KYPuFE5XaIswGNdy7Gln5ibuDieN6/6YLGJ2h3d8yS
Gy/1CvbkfhIJaIPC11JFCEWFrcGo78rqdTk56/PGgFBErqrRWguLLMviEzmaZhjHmYtJ4KB8mZWY+vKHNLPrqyg+vrW9xFhmrvHetGFVZI6ydLdSYo4lxmqA0SE2F8pk
Qw3g9I9xQ3lRpTdaraWrWvFbHPbxbWfVxXkqhmZEvxIqCEz4FovFchLkdah9k6RHU6bgO2hzpVM70iDAxRsbW8DI4k6l/Kxkpzgccw97EH+STKcYjofvHyr6qf2GdtEn
PalSfV/NFJBjz49Sizhk9+ciDPTnZZazCr2nLu1ibwvhc3JgWOXi63hzXHJASXLAFo18HxmdTOboTvhkhU63iDKVI40OtFdp15GOTDduO5GaBgmuZEkASg5OzfQecgXm
BM+zh+zUAfEtGxg+YznVe0e1Z99X9r+dAMMtGfkok5RHOQ+GLILdxlsgLvYveXE7IlBtUuRC4KyvcV0UaCUqfEMN4PSPcUN5UaU3Wq2lq1ryJGO+rSjRl3AeuzqsNGyF
62KdYBvglCTslv4sBKu5LdHlKFEiX3hS8GwLUzkUmcnACl1+twpO/o+5Mel8eysdeIRzXRNIEzQvj18azTN0UiwG7KTeQt6KNMpS6FCAbeNDlb7zYMS1+i3p5EHsBLLY
bR0ky6XrOB4czEonuEuRisdQU9VStljaPzTQzHKOJXSh0fXnAqpTWGV3UJV+6gMNlM9LFDk5XemfePQjdp0FiN/KBIO6Bqayd4mKcoGtyo4fOq4ypG/J4ISgKU14U3kM
WLEltZ/nKkvHzJEhgE1BiuEVeYBtHot7eYFbO3lBiAFLNYsurzwS5IIyc1uTOM5xv5ULOlt8QBoVft1iP22YZvhg4uFpjxHx+eQZNNg0OvasMK61Cvgg90lJy8jCVQFD
961Kjjok0iHYUyDIOR1Yrpz/RZyy9LJlTGCOBh5y0tlBd3zuCKbj0ZGQX+Q64sNV5yIM9OdllrMKvacu7WJvC4k3CDCL7eg2pAm0gAq7NcZcoyyP0oBmJRjbQ7yYAE0w
zSU+SAcAXhiVU6sk91xVrsBOcKRSNrPco1YF5pwPwV8hx+FRT2g3+5VLtjyyIr6ZlM9LFDk5XemfePQjdp0FiN/KBIO6Bqayd4mKcoGtyo4fOq4ypG/J4ISgKU14U3kM
WLEltZ/nKkvHzJEhgE1BiuEVeYBtHot7eYFbO3lBiAFLNYsurzwS5IIyc1uTOM5xv5ULOlt8QBoVft1iP22YZkXn4NfdV6FGZpAyw6JElIdyn0EB7W1neic2RU7pUpJb
U6bgO2hzpVM70iDAxRsbW8UpV4/EkMTFdHjLeZsJFAjV6kkvwL8hD7Qtuy2VqP1DpC2WC+rken9jA5fw0Tn6eTNybndMlT0i6KDi8fGbkHvUjtq8y2CvINBje8Yenfas
spgc1EbAyNk0QfeJEmgDV3MFH0BnTQ6X+8Qe88VOpbLI/k+T/HYul4nngNWCZd368PUZrvwHxt2PNViA2nWv2hXeB59sqVE+vBU3J2zNCaOkU6INqtNgQeas/q9Jh2oL
Ym7g4njev+mCxidod3fMkrSzYJ7twH+f2N7yX/fLbCJFha3BqO/K6nU5OevzxoBQRK6q0VoLiyzL4hM5mmYYx7+XueWv+aVxqYz7x5bYBR5yn0EB7W1neic2RU7pUpJb
U6bgO2hzpVM70iDAxRsbW4bDm0aq9neYJwLi4mTs2h8MQfBqD8cEHq2t4g6y2hRwOewmvw0BJZCbraGnzYe4daw4HGns5yTPlrVLa51nHdw0kdaLOix2tEuYezhKONNt
Atz0s6B7ERBlT3wsmLyw5NHlKFEiX3hS8GwLUzkUmcn+lIcygWeWN0HzpKuXevNlAscK1qwacUNjy9iaqL7kaLOtjYKeg6I3dA6oAZkeB9qApAx3UF2iCArPHry/wIYr
UwZqFrmctMiWvohlxEGfRWMvbolzBbggIGu7eVk/zGltTScrpZfW1JT1UdbngFFpLDjBiVxeQUq0Y2n9Z5lyMEURzy1m2KMx2qi1KpLRG85i8PBDjUU4gilcEz9ZWSaV
bHvgagnI71cSObPvvIu44amtAxvBqmFlO0ATy8GPLY6ydLdSYo4lxmqA0SE2F8pki/7P8e7ESyfLyrpYbp24Ym0b57EhgNiXR7bL77f+CqzR5ShRIl94UvBsC1M5FJnJ
/pSHMoFnljdB86Srl3rzZX/brzwY2Y1tPzDAzGZyEju5NiGEJoqDq716e+XXtHYDMyn+ub6mbQpqFl/WaNPKrWx74GoJyO9XEjmz77yLuOF+y+WsZ5PSoOqT/YHCIm1J
0Xe48InjjfkmxcrQJbF7nipaZ7UDzn7J6YIE50MMnSpJb00XoIoG4ct2t9nx0Sr2L7Eqynp8XQdwhfJZmFHvTkHQQdD1O/BFa+56rVchl+2cE9vAwbaLesFO1z9QXA5D
jriEUaKCbNLG/fe/9dtJlf7jpIisLIAD8dNI5F/3MBf6WoesTmZS/vLduoF2M0FcKjSSNhGh9eaWp2daon/nCZL5oQj7lUrrZ0XKnjXlSOtkx/BKJOOGTBa/SaAH4ckJ
ev/AYIG78lNWhsflAMIiZtSO2rzLYK8g0GN7xh6d9qxJIpVN9ZhWTh3Gu6+qg9ApcJ3vhLd9TxAfhiA7i82U6BbeAHwPJn4oV8Fr3zbpYNg+jYQ1+aFi9BI6UFxAY03L
yijZh8LmwfiKibX/WkCyZG/bD9Of8txvgB7S2FMwos9QO6P0Ffi5bhAiJhKTLw++eWKIFJaYwMT3ip4k2OqUHRzcrv/vsQ03RRdpYvi5bV9EVzjnqYHqyYO0JtwGVq58
VjYYvNlhPzr0PoHUOztllGyoExnkgn26/Crp+Tkkn5Px/Q5G1LxDqfQyUhrzX9fgqC8FN8TpnE/kVLIpmNKkJSr5MAewiYKHyGuBZXk2xWU9gMj0oDKltzdQmc/1krVB
2/bKtlshAIdjfLyduhFtRp/ntXmEZs8SNiAVj7UC6+YyvQ1z0lbgYH1o0CmLcgaLkDW9c7+okh/55lO9SPVExgtARHUIwtZZvOJpfyXMjeiAS4Bxbh2FZhj5WZV2bRJN
C+w4FNO3uX7hTuNOMr163mmf2aei7L5Xm+CDjTQOb4IW8L9zKzQ3ZeLeMA9SnAUKgMjrZpglksZBGY2K2V0OkBC3sUcqk0X4YVBAc1stI7YCrKWwkulLNin5DOn9ebhX
YcQchLPymHl17LByH814+lMArvqfdj1OM1u4OuwLpvpXGkEJGnb5uyM4rmsS/WDSmgYJrmRJAEoOTs30HnIF5nWP66LeE/IObZ1MiQBqT4oSkteL8YU1X6YyuF8LmUbW
jDErLOIMfzrmpMUoIU8meCyREanivoQCwP7zkgRIWbZibuDieN6/6YLGJ2h3d8ySK98tpaXst3Ly6+u8y+hYF0WFrcGo78rqdTk56/PGgFBMADb3QNU+6p8eFD3nXm2v
UDuj9BX4uW4QIiYSky8PvhFpSNYdg1SLxSOFREyYIkulsUN6hfm/tXNpZmTH7kybyijZh8LmwfiKibX/WkCyZAwokXyLKmuwoSV37jr2myAbP6mdLE3iq8NKmw32NMjE
b9bIlrN0iF4ojiVJUCRBxBaNfB8ZnUzm6E74ZIVOt4gylSONDrRXadeRjkw3bjuRmgYJrmRJAEoOTs30HnIF5ndf3W4tS9jkUXMB141eH4RB0EHQ9TvwRWvueq1XIZft
L4sq+aAK2V7ou8drubJ8BJO+lCBL7wwwTR+vMtdngtmUYHUA9G2m39fE8UjAohUl9vuus5H+VJNn+frGjkcW7qmtAxvBqmFlO0ATy8GPLY7ZuhdCSW8d+uW5dgM6Gxcs
w1TuIVAwx/S2E+hhdQqcjaHR9ecCqlNYZXdQlX7qAw1jULoFZVG2phyu+RZn9qpc1IQeVeng8oIPPdg3BkT87DvmDRagm2rhwFKp8j9qtv8fx+He3AxyLmudYrf2T9id
PMVdP3/wwep7+Z6U/kKzzvX4+JDB1lGmzlJaLYpjjJQHjthDfcEUnWy+SAP9bwUi/lk5yq2yHCj/T43XG8QCtjwGN4HX9N4tLE4tFYBfCfXtXExFVPfwxcfPB478F5DI
8FRbI5AVt/OKBT3X0EKIQ0xh2EBT7q7izBqrDhJHWq0jk6S7sFr4XxYBfWAPfJXSXvtM1nwaoXKRxvOjwm6lCOp6TppMZZELsjOxkAwK7B7ZN8lZfCnffRa77vzwM0Nd
RVzxX2djx8nzqhTzJF2A1/GMbgA4zugJrfWQXfsuV1yPQzUtl8K1qaJ/I2lvNr55SOAn14NbDMj38+H+j5B6TVp4yWt1Id0LlEuhiACHe/4lmH5qmvoRCwnUvU1gfW5A
+R16l9ZUHhUdoU8nS1FVt2xSMYBkuy3tx4C7OZz7ES+wahFXBTWb/mxWQYhcD6lXdrD/1LQEYqFUArU5KCN35yuIWjCi3WPbKkVGHNBR5fA7iDj3d1b9RYyASikdDf/2
Df6PEbRqnNmOORAx2eSxq3hRWBBzrmYuy+mv7t7zxs1VjZkCbUig6Xln74dUqo/wzpENFUNkSyKV/XC8/3+rvNexkOUXK6cHQ46W1ypRN27sbqZRQH8wcNmDgsOQ4AUo
vcmrvRMafdgjCSHEQGkd3S/LdUT8ScN5tet7zALclV8lnnR5y1uVy8F3I3vJF+z9kf6xnueXRW29OahY9ctBfEkJ9FIU8NUnXU5IsaP8mhe1r8PqA/G/wMz2IhMDm3vk
BWM66DX8cyPJZiGnRxdrZ/LXidYVbyT3A7ftdlFkytajPR7tKWRB+Qkz91wS0VpTbFhGQ3iK1IUreSkhRuLCRm8ps54CzFuooI5/gjM53nNxnHU1NwDkU9VhzNnVZ1CY
764KGnKnKmqsv7O2E8G182nKugTY3CZIBPFDeJHfFk936BBwKC1+kLAQZ9KHi6BYTJIpufQVZ8S2+uTHNqgiqXl6yzhVLlcXtxiohkB0h/OlXMbVF2Sf2yuj4kF/3wAV
6E3vYQQKJcZ8RFZoT2XkDkSH3Yn2NXSoS97obiyRD8X1+PiQwdZRps5SWi2KY4yU3AeB1W9Td7vCUHEKBQ3RFv5ZOcqtshwo/0+N1xvEArYfv8lKki1LEC874PZXUy9g
7VxMRVT38MXHzweO/BeQyPBUWyOQFbfzigU919BCiENMYdhAU+6u4swaqw4SR1qtZoezolv/M88CeyxkDlZJvV77TNZ8GqFykcbzo8JupQiEuIKqhzWxQcQf8kojazTP
2TfJWXwp330Wu+788DNDXUVc8V9nY8fJ86oU8yRdgNfxjG4AOM7oCa31kF37LldcHuAJSq9YsOl44Fo6CcoO40HxVES1KPMBfMOjWbqllSL1+PiQwdZRps5SWi2KY4yU
/SQC/MtsLMmvaZJmw0cJ8A3+jxG0apzZjjkQMdnksat4UVgQc65mLsvpr+7e88bNR3rZlpqk7GqZRBIsRJIssDhk7HnIIH2FKV0CR1LTaG/xjG4AOM7oCa31kF37Lldc
c6D8Wc3SR4ftd6hjfov0mAVjOug1/HMjyWYhp0cXa2fy14nWFW8k9wO37XZRZMrWyTJFMFuw8+mEg25bjmgnxoJ9palBHxB7J/vAPiRLJQp4UVgQc65mLsvpr+7e88bN
A9vNIZVHzeWkwuFpKkwo3uhN72EECiXGfERWaE9l5A5Eh92J9jV0qEve6G4skQ/FLiu1/onR3hqI8hH6bGBVXdntEzK/uVAPuKqqRjJ95zPmzEsNxKNVcJmT1KY3NJQX
DzVic394AG5p5fa6URmQjWEGG55t5AbQMJ59PA6B1DUrAPdNEv0tHaJWmhljYdMxBKTYJ2IFZM9Ww9TNuK3ozDcbLDualpUjeXbhRhsXBuXAwr16kqVYAYPBmuHDF09O
QzZdyyA78q9y1xAqWK00fjmpCKliKcH3ufofDcqKmVnGJ5wXctGbYmz8Iq0GzWrZklLusCDtCsdOBSjoV/EBqd9LY5SnKIrKZT6HeYdgDkrARNxDjvnTawzfBXZgYA3t
3fyoj1p1pmJtZj99Y8TzkC81q02U8t8puUXYClLzoTdMXgVoJRb4W2yqfWAf1COiIRiWcKa72d76UaFxS2fsLFpYq9BpmDBMZVJVPqkyxIPrDG6km/r/scn1Y5P6cq35
jsXa3AGW4NSr8o4BYK/fJxrXH90LEW5y+xiFYbsTprZeix71AYESwtgJyC6+yG1BRDTKJpdEx3jv5eKGVJmOCjDT+QHE53wMFka0n3eM9DR8Afp+XuyDitLK0QlQl0CR
LWPVVTOxK2/flPzy3L518zDT+QHE53wMFka0n3eM9DRHnlhWbh8BgKLaL77bmdgJEyZr0o+ag4BMdPN9QWdW7zDT+QHE53wMFka0n3eM9DRMfuKKPbmOCKtiOHmfrcyK
i+ema7Mwkdj2siSVkMArVDDT+QHE53wMFka0n3eM9DSXH35Kac1qy+Gbpj08ac7Pf/OzYpTJn5sAxW4d9ci7h5ARoxAOYkatQ/W7azAhVaZGIeLuMqvRv2h7xH7ld2E3
ntyK8YmWZJEk3wlFTp17OZARoxAOYkatQ/W7azAhVaZ8Afp+XuyDitLK0QlQl0CRcC9i09bXQ1enB7VMtlEDKTDWTaUyAvX+UdtO+yuW/LNf0JA1ypW4RKCIrdTCYr66
RH3313SbhY7b2rkU3inZWu1cTEVU9/DFx88HjvwXkMj5eAiLDJo9akoIwtvYnM4dtlX4wP0wqLOx2FM40e1Wc8BIyc0Pr4LqCe2iAXxEhgJ5T+7wRuMgejgAtEorEicW
dGZUh9kt+Y0zoRoAO6yo3yEAix6j9XVISLooL4dOW6vDw3m14bxdFgEQ5cyrGRiklHulFGq+aVjS157D1XJiO/WHpsqIfbOv/VKCtqwcMgL3rUqOOiTSIdhTIMg5HViu
nA1FNaOg4Awq2h5IPHFYqL12qNT9nAHC0Pgx/KpZP7KGv8yIEHYrNmT6oT3xp/LS/ArxS/Z166l2bwIqCG9P+/YbHM9hBaNjUxq7HTJJap4dooeoAJxYmBCwQRH4Mh5S
qk/vXKTCiScx2XksuatAsFp4yWt1Id0LlEuhiACHe/7dJFcvwReiZgZFyk+WA8Gi+R16l9ZUHhUdoU8nS1FVt+v1mK1Kgwz25HiWwPC7RqCdG77qT0pL/25BPXQ9DqBy
RqTlt6pDI4CejELhPJi4ugyWIeZ1q2mW92I6Kqo/RpUOGn7G8Ah967tJFli7Gi+r4RV5gG0ei3t5gVs7eUGIAUvgi6gwoTsxThHs9gfVe5yR/rGe55dFbb05qFj1y0F8
aSyy+cxJn9/TUbFVtMjA9HtRUL2lelZc55mZLAI6V0myaFsLREpynj3bBx7tCjV7CjSwoDtLzBPOS5hvItIQlw3FO4TsMI7oEWyADwwxjAGFpTkeJHeyQGzsX4DaHyZ2
oCir7M1nfcHuZU1nV6UOvr4t7PnkBQyUjNxo6manzgMBJpQFvYSo5IpgUGHcU2dYWOxC5Vtj6gZM17vPVRtATY7rQlxX+xpmWJBpiBzCG1uCfaWpQR8Qeyf7wD4kSyUK
cxhWf0TB/upgCU06bZiwUlWThAVyFv05K3WNK/oN8+WLmhX1swEDi4ZrfgrTW08QBWM66DX8cyPJZiGnRxdrZxRUEz6Klq41wQ8/83Yo1g5vBYqUswwx+FJfjznPGfs2
hyTYnOL+UtVKhpDI5GCyrUd2PBkNf5YWwxKad/PFFAvvrgoacqcqaqy/s7YTwbXzdhQMM9a7idBSSE8qGgdhacRR260H6Ind4S6jwUiojpAPLsk0a7laQOH33aVInT84
/8qpbMLyB4E5VoP6KnLMD0UGAmTmNuMp5uxmQGAh4WBVjZkCbUig6Xln74dUqo/wvsEMia04GMSi/ypp8l6XIkLy8T9m2pSXEImNNbgcHtNGQXA1sFSXzrOuY1sEsjwK
4Fp6WJo74ahkX1EQe0WyzAexj7Dhc+zupig7gqNVkEZCE0zpOm9TIegNIU1KHwM4hOqDpXeLEZ6xH2RJn25q9KWzxny7Ra+XM6Xoc/jzwWxhGfOoECrSy+Pu4CKF8ktL
NXkewmH8Afa2dQGaI5KFadK9yhVK6bl7w0BLKcRLg9Bsxk11mtRRafkcMAKks1gM7VxMRVT38MXHzweO/BeQyHG1mRLLIV1w4iBgW4bnER8hTWydodF9eFS4+gkt08HE
AcTvF8gwooMKmKArv5m08HNuLEOg257HPV3Cz45hRWHZN8lZfCnffRa77vzwM0NdHAjSM/scI0tUO+Dvsn3uvOhdtTRBIr0YN4IFF6600+5Yxi3NlPexomBxvnpsgcmN
523Kd8J26iNO41z0v9Tb0hlyV5xaclzhtXTaXYxgaS+erQzZxXX2JTV/LGGbCY72vXao1P2cAcLQ+DH8qlk/ssJQCl23S4CcLj8ixtv/ycjyUJS2vOGdYyNCEK1cG4fW
s+rOB76DbYGn50lpAm8GwMav1Hqb79sfMnPXXpb1WZzOVe6QjbM1C5NxkJCBGWmcjj9T/qesR6d+TD5bG+PaKlzzsg5NyAtJpOhm36VgeNSlXMbVF2Sf2yuj4kF/3wAV
yWIGw/ij86CT2VvbhU8N9lrelGspI9p6l8CDq/Q/d0qLyDxeAxV63PfuxoqmECOJ2P2YUSewiuiDFKSrzglKEA3+jxG0apzZjjkQMdnksasgPXHZelW1PSuKe6FILjm9
eraMep6T5+iQeNZY9KMyuxlvc5z4G+9WmRekXDSiIKt3rhjws/ZNPBiAsDEBq3+kvcmrvRMafdgjCSHEQGkd3TG/wNWQk6OoIWb8wsvwZobLMaE5OyVxqCFRwfhjLQ6X
bFhGQ3iK1IUreSkhRuLCRpjDvRbJns/L+ToJWVSvpo62VfjA/TCos7HYUzjR7VZziTD+rF0MQBTYCFAWi+uXOwEmlAW9hKjkimBQYdxTZ1jKxoniKMra8fEb6gh1ndKV
3TiPIjYIzHEcMVbOT+Ff1BFjzToxW7vcXsiEx8kE6TyfuIwrTKm1hH71b3h2shrP7MuvNyT/ns7/0Qr+G4kJnrX0ef2dvipUg7MQGSQt1L1aeMlrdSHdC5RLoYgAh3v+
YhoPvhA5wdEh1U+YMS2li0L94zviHydJ99mvNKtQZOcmgi/MMqOCI7U+11cjUP7tRLrlFGzGbU8pwLxt+j1YoO+uChpypypqrL+zthPBtfNM6R8T0XDY6/WqWXBqLMrQ
IcPg8Ps3+rTu+CiXszLrA50kqlcPP8B6kqJ8iwPf7FhjXJyz/PAtnaInCvKoMz5nQhNM6TpvUyHoDSFNSh8DOITqg6V3ixGesR9kSZ9uavSls8Z8u0WvlzOl6HP488Fs
HPWPKmmS1xvXkoKfZ9vvxXlP7vBG4yB6OAC0SisSJxZKCoZsenvf8LSeK3rixQeKdt9eZ+f1zYVJh7b8MzG9Rr12qNT9nAHC0Pgx/KpZP7LCUApdt0uAnC4/Isbb/8nI
GTB/IhiL8Uy/fVV4+ZeeOZ0bvupPSkv/bkE9dD0OoHJGpOW3qkMjgJ6MQuE8mLi6iKCt+7KYWUuq2+n8OvIdlwo0sKA7S8wTzkuYbyLSEJeqMmpjIPJKd5qVJdjgcpX+
W008aip6jOcJ7bL3jTPBwmxYRkN4itSFK3kpIUbiwkYGvKd5xD9GCkG6DscErtedVZOEBXIW/TkrdY0r+g3z5fZqQhedztZ6TqOcjZSifKLsy683JP+ezv/RCv4biQme
yGMwB7a1f3x09oFvB28mp4eaAN5FP+c4Kp6PkO43XVSdJKpXDz/AepKifIsD3+xYO4HuAsPEbfOA8ICfnWazEkITTOk6b1Mh6A0hTUofAziE6oOld4sRnrEfZEmfbmr0
pbPGfLtFr5czpehz+PPBbC062GUW+EsEA02j1CoKIpt5T+7wRuMgejgAtEorEicWADgxkC8TTlggSOQLSUnqW4uAwo5CNwJWmEZRzPPY+7u9dqjU/ZwBwtD4MfyqWT+y
wlAKXbdLgJwuPyLG2//JyD+sSgp90/Wew0n7PFopsOqdG77qT0pL/25BPXQ9DqBy48tMwLZuIDE2TSZaZWh4e03qGBp/YFFnNgW3xvAgRecnu8ZBYr3GwwiJDls8bZWO
krkW/f0YUNpaDdURneCMr0cNJY14ITNjGEGaIwgExXF3zF62haLu5LbsbASCEwYOyLcP+WhkY5XAff224JTIk5ZvQoINFXxyi0Hyq3999G+VhXH0DhPx3pryBuATixQ7
+fxcUWeEVkYFn/b2sVnL6EHxVES1KPMBfMOjWbqllSKOMFDvk8QYIBnLjEBA8+5nFOE4RApn0hcntkAaARytsT9nmw7QNoGEmwXzH6I7gflc87IOTcgLSaToZt+lYHjU
i8g8XgMVetz37saKphAjiWwH0K+yxpcq5Y00V5MkSvpFeUvL8R9oXQ9mAwaXACmyR59trVvR9fbyKqNIeffW6o4wUO+TxBggGcuMQEDz7mf1lHkShXjS02lCFn9zbqdP
/xKVZtreaQx/tCmlzC6KXSXRJHovD7IAenFpPBfPiMyCfaWpQR8Qeyf7wD4kSyUKeFFYEHOuZi7L6a/u3vPGzZoiPd+tizCzzWWfZtpSw0Y1jXbnNUg0qKYldkDMMeg9
2Jur6G7mh/IsPxRFzCGbssqIJtEmvYeBjKtfeWMCbYi2FzhO9lN2Qa475Kjb3Bv+OGTsecggfYUpXQJHUtNob3R4VmpRttNch5ggYOmlF3b3rUqOOiTSIdhTIMg5HViu
fhiMltqcp9Dx6Mg2MCPw8JZvQoINFXxyi0Hyq3999G+VhXH0DhPx3pryBuATixQ7IS+x/MSxqpsQ7mLPhZ4YWEHxVES1KPMBfMOjWbqllSKOMFDvk8QYIBnLjEBA8+5n
FOE4RApn0hcntkAaARytsVO8n3GE7Ywi7ibUXf/Q3ZFc87IOTcgLSaToZt+lYHjUi8g8XgMVetz37saKphAjiUXGLoSgA/CfSmQ7HFWtGmpFeUvL8R9oXQ9mAwaXACmy
R59trVvR9fbyKqNIeffW6o4wUO+TxBggGcuMQEDz7mdj/pJyKo+8jX/gmT948Yr+/xKVZtreaQx/tCmlzC6KXTvvlU/ZDu90xhOJabtjz1WCfaWpQR8Qeyf7wD4kSyUK
eFFYEHOuZi7L6a/u3vPGzZoiPd+tizCzzWWfZtpSw0Y1jXbnNUg0qKYldkDMMeg9TCH2dhdy3Zj7I36Sk0/YRsqIJtEmvYeBjKtfeWMCbYilXMbVF2Sf2yuj4kF/3wAV
OGTsecggfYUpXQJHUtNob3R4VmpRttNch5ggYOmlF3b3rUqOOiTSIdhTIMg5HViuUgA3+YTk6QnAIvqpnK8sj5ZvQoINFXxyi0Hyq3999G+VhXH0DhPx3pryBuATixQ7
/aGo3Pp2MuK/2Bi20P8AVkHxVES1KPMBfMOjWbqllSKOMFDvk8QYIBnLjEBA8+5nFOE4RApn0hcntkAaARytsbd7mS2OjUW8JbmnNDSH2oVc87IOTcgLSaToZt+lYHjU
i8g8XgMVetz37saKphAjiZZqywg8HtYkiI02Q6MktKtFeUvL8R9oXQ9mAwaXACmyR59trVvR9fbyKqNIeffW6o4wUO+TxBggGcuMQEDz7mdiUYOmBxzRsHI2yMihA8yO
/xKVZtreaQx/tCmlzC6KXXbfXmfn9c2FSYe2/DMxvUZMkim59BVnxLb65Mc2qCKpeXrLOFUuVxe3GKiGQHSH84vv+0sdQ9IRSSIe0MBUl3tlQIBpSeXvuEcpZItP2pDk
LsPkAvDnFNce+xq48VVa4cqIJtEmvYeBjKtfeWMCbYgwd2SXNxJTQLarsfdYHtvehQ0RNiV35S8I+2BGyV7tMxN2et1M5Ga441dH6MyHpFqz6s4HvoNtgafnSWkCbwbA
7g7/hSrYDjzhNs7vGgMIJK4DbVOFYVll+TcqGEEqSovKiCbRJr2HgYyrX3ljAm2IM3Gmks5M5haqxBIqacsYIc6RDRVDZEsilf1wvP9/q7wlALfx/UklBgBv0bODmdcw
AcTvF8gwooMKmKArv5m08GzKhnWgyxWKSXh89+FjSZ3wmhKcAdZpTC5JXOfkY/oknRu+6k9KS/9uQT10PQ6gcsuva42DkVw9fAapLLIvv22dG77qT0pL/25BPXQ9DqBy
48tMwLZuIDE2TSZaZWh4e4AI0oMGi6KSjqf7m7DGyu1d3h3L3+RZPDXm+Iy9vJvuzlTj1nIAuz7guo0S0NkJZLlGp9GyyVXUIl39YNIkwOOIwrL6MXLjcUZecYFvqOnN
FcGn5J1SJmuIXjcwx1okEhcg+fBD4uS1oa+3MeajEqf8CvFL9nXrqXZvAioIb0/7WnjJa3Uh3QuUS6GIAId7/hcOzWn7t9K9LES96qdJZT75HXqX1lQeFR2hTydLUVW3
E3Z63UzkZrjjV0fozIekWrPqzge+g22Bp+dJaQJvBsCsJE6/UkA5tB0aQGmDMFiecGtOv1mIfOD0+hN14ZsB1sqIJtEmvYeBjKtfeWMCbYj2GxzPYQWjY1Maux0ySWqe
764KGnKnKmqsv7O2E8G182nKugTY3CZIBPFDeJHfFk/xMwnCSwDOdR7CjlJLSyEjeXXSW6XSGLk63+hr6EA4cn86EXR9e3+KE0EmfFCGwej8CvFL9nXrqXZvAioIb0/7
WnjJa3Uh3QuUS6GIAId7/iWYfmqa+hELCdS9TWB9bkD5HXqX1lQeFR2hTydLUVW3E3Z63UzkZrjjV0fozIekWrPqzge+g22Bp+dJaQJvBsDuDv+FKtgOPOE2zu8aAwgk
c77TXVikYrXHqGwVzZ0xWMqIJtEmvYeBjKtfeWMCbYhGVqqi04rYuRFgncgXmBBw764KGnKnKmqsv7O2E8G182nKugTY3CZIBPFDeJHfFk/xMwnCSwDOdR7CjlJLSyEj
eXXSW6XSGLk63+hr6EA4cujY6DB+cIprgvHt7i8WCH78CvFL9nXrqXZvAioIb0/7WnjJa3Uh3QuUS6GIAId7/hflEgB9zcQa2NknP78o8hz5HXqX1lQeFR2hTydLUVW3
E3Z63UzkZrjjV0fozIekWrPqzge+g22Bp+dJaQJvBsDuDv+FKtgOPOE2zu8aAwgkau5KKQnUI87HRHRcOVgxpMqIJtEmvYeBjKtfeWMCbYj3U++Xx6DXEPQuk1JqWKgG
764KGnKnKmqsv7O2E8G182nKugTY3CZIBPFDeJHfFk/xMwnCSwDOdR7CjlJLSyEjeXXSW6XSGLk63+hr6EA4cuyF9pJkSjio2pp7u5qZXjj8CvFL9nXrqXZvAioIb0/7
WnjJa3Uh3QuUS6GIAId7/rY+rdNDrivbm0JWn85G4E75HXqX1lQeFR2hTydLUVW3E3Z63UzkZrjjV0fozIekWrPqzge+g22Bp+dJaQJvBsCsJE6/UkA5tB0aQGmDMFie
uiqhS3pL+5zF4BwJqHYYTcqIJtEmvYeBjKtfeWMCbYjPU0n/37fNjZSMYUxW5kLb764KGnKnKmqsv7O2E8G182nKugTY3CZIBPFDeJHfFk/xMwnCSwDOdR7CjlJLSyEj
eXXSW6XSGLk63+hr6EA4cjQeXhUGMjfFLAaxlnBjiCb8CvFL9nXrqXZvAioIb0/7WnjJa3Uh3QuUS6GIAId7/jcoIblGrtAbQOUl3uCaauH5HXqX1lQeFR2hTydLUVW3
E3Z63UzkZrjjV0fozIekWrPqzge+g22Bp+dJaQJvBsCsJE6/UkA5tB0aQGmDMFieNYrlVu38x52cNDiWM0s+m8qIJtEmvYeBjKtfeWMCbYhEuuUUbMZtTynAvG36PVig
764KGnKnKmqsv7O2E8G182nKugTY3CZIBPFDeJHfFk/xMwnCSwDOdR7CjlJLSyEjeXXSW6XSGLk63+hr6EA4couYq4zXBcsMx0KDpzic4+v8CvFL9nXrqXZvAioIb0/7
WnjJa3Uh3QuUS6GIAId7/kQvX0Tu16L69Z+/G1n3O2wwGVsPHWOurJQ9IarTTx0qbymzngLMW6igjn+CMznec50bvupPSkv/bkE9dD0OoHIRpJnZ/fOLDOSakT9ZoPoJ
fjG/PhBai45h21hbDN9fmMqIJtEmvYeBjKtfeWMCbYhHetmWmqTsaplEEixEkiyw6E3vYQQKJcZ8RFZoT2XkDkSH3Yn2NXSoS97obiyRD8WOMFDvk8QYIBnLjEBA8+5n
FOE4RApn0hcntkAaARytsRGmSG1aByIIbLuarGdxoBZc87IOTcgLSaToZt+lYHjUi8g8XgMVetz37saKphAjif5KjftS+Jg2TvZENZAJ00EKNLCgO0vME85LmG8i0hCX
eXrLOFUuVxe3GKiGQHSH84vv+0sdQ9IRSSIe0MBUl3tFB5mCG+9vO2jZBabC85SdwHFAE0RL9TQ5ZspaHCNkB/YOXjc2w1gU6tZCQaytV0oZKadloSmWDBChbLy7Sskv
BwYK2HiqvYtmyzGPxj7Wdp+huwmO2CEdblV3OUBp+Y09pX1b1wM2ldS7tLU3i+rFFbzTlAgNdxmA8Eb65WjIqplI4A8ojStoMzDETEuUux2oxZl264ujB7TBmJ/Nsj86
/xKVZtreaQx/tCmlzC6KXVByGZP2k+AKzoiCUlBkiZjQVAKRbKE2SmEa+qd/YO7iyogm0Sa9h4GMq195YwJtiN8grni+GhFq4bTTMr5bKX7b34VnHE7vFMukW0S2HoW4
J1FSVRlk1+4Vs6GZYtIgRYvv+0sdQ9IRSSIe0MBUl3uL7/tLHUPSEUkiHtDAVJd7IHg180fdhXf+klUV/k8q85n+mNwrQORPk7mYkI/FboB+Mb8+EFqLjmHbWFsM31+Y
miI9362LMLPNZZ9m2lLDRmbA16q2uFZV6MOpQP9aD6xxQVnaDR5XaZ4sfQI3j500uiqhS3pL+5zF4BwJqHYYTYMBMgC4+wYeG/dpQmR45IKFCOC3bn5fY8EOkW5anCmJ
Gn15UcAfq6u0+U/spP1dn+PYpK9igx5sBhjqKI3uvc8yXGTO3/azth3u1cxfk9fav7f46UcmIiEjRwuSxqUWXswbnnRofqxYq0XxNb4cb3EBxO8XyDCigwqYoCu/mbTw
AcTvF8gwooMKmKArv5m08IoXWrSN+MhWs18kdnblMlkqXJlyes5xjMu2lmUDTqG+WKIz9Q9vwx4R442Tc3bJrxXFdsdoz94eHkH/bkJZeUcKx5nfTZ9ni8au/H5bvlVH
c8HatquM0JhWYhr6G8/iGlzzsg5NyAtJpOhm36VgeNSfhuOVGSk5et8oamBA0TsiEORVO6rfy0QQJf9MTI1bevwK8Uv2deupdm8CKghvT/uILrfrHIjBZMi/CWXY5LwB
zv5ocQ5w78VGfgs2/okcIwoy8UFCPYIs6jh56ks1zrX2Dl43NsNYFOrWQkGsrVdKGSmnZaEplgwQoWy8u0rJL2/wrRUdgqGbghg9XXcFAj4xZ/ZbSNQRh+emJiIW2GNm
ysVVXUEulep3m4FXjNsuFH9V5lnijLjFn4O8rkIRQ2RwmR93LGumvYHQCwPZIxoGqecQ7dAdIMX9tVKdzeuh13j0xHZrGynF19sHFafYSdjKiCbRJr2HgYyrX3ljAm2I
FyAMhSREoVWGAOzEl8PBRjsnlJ/1dG4tJc5z0KSqbDvKiCbRJr2HgYyrX3ljAm2IPqW6IxEbjKdi2mssoy2N56P/9KuXnvdZV/2sQdsYs9YGix0rTNlai81EvHiJC/ec
nRu+6k9KS/9uQT10PQ6gcp0bvupPSkv/bkE9dD0OoHJTox7uKKy9nch7O4kKWSTDn9d18K6lIoFhW0QCnCIkw9KcRz49trRooAAcgWslHwqz6s4HvoNtgafnSWkCbwbA
HlBzl586tzQeUagl27WfRgaWA51WGjoGfE/k+bY4EPJsSlZVR+Hg1tQIdUf7wmDuZru8lh/MIOUP49cxjApzNwLqmmD/XRgzROTTtk8GkUAmKSWLDdKZsgRUqikO/M26
HmcEzAtP6wSVwuUCrOrzcHyS/X1hroLe2goGfk44QjUnydMvfwRZAv+TdeBxYytSWxl1AC108omuYnUm2r/X76D3o7lk2075mvR49GFcOemg96O5ZNtO+Zr0ePRhXDnp
CiXztXH6JOajxg00z2JzOBmopROpNqZyDZH/ROt+h5/b9sq2WyEAh2N8vJ26EW1GFOE4RApn0hcntkAaARytsTYGKzF/POZMdaywOU4JFeHV57rqAx6J9vL4DdiRROPN
/ArxS/Z166l2bwIqCG9P++PLTMC2biAxNk0mWmVoeHu1gJN5rZkM0bjAOJLgKLTk/xKVZtreaQx/tCmlzC6KXXPdwrHamSzKYG0wNeo+Um9l7pAYroftzLbLO4S42s4k
/Mu4YceT9gf+atJJuVAL+PG9Kqkoxg4HFe+4g8ZlLHTxvSqpKMYOBxXvuIPGZSx0N4oJEtinp7R5kaF6yHBAggPq9he/KfROBeef8+TQxs9kkKgh8rvzI/x6eVVPEPSP
/wCw8Z9KwwNpYlpQeXe/vyvQL7JwuseDYb+STQzncqS6jXT/B9mLkHW0G4MUKPfnTCH2dhdy3Zj7I36Sk0/YRs69D6VBaxhyBCpZ9P1MhBugim2aSZjwmakm4rOhr9L9
F/VqdZERRiQuDgNNqud7MMqIJtEmvYeBjKtfeWMCbYgTLBG5dkvp3OWftmBxTWC5bnXe7P5GsdRsJgUs7swkP5oR3q48SsCpDd1ryOxwFHVibuDieN6/6YLGJ2h3d8yS
Ym7g4njev+mCxidod3fMklPOyxMOaLh48ZgSfBQx024ND1aqudAbBhjMAzWHs3YJm7OUpyqr9qjffPe27Ox6AvetSo46JNIh2FMgyDkdWK6OfyoitHTO23+3q4HrZ2re
sg6vlhsSUprb4u8exFX93fCaEpwB1mlMLklc5+Rj+iQgcPcbUsx1O8jsW9itWtj8w82dHOCIJD15TRF9PdWO41zzsg5NyAtJpOhm36VgeNRVxGkaXeFE1f7231cp+vlZ
SiYo+yKduN16M+dLhgqK7Y4RTYa0nyg/angvDZqKh9DKiCbRJr2HgYyrX3ljAm2IYqtMmuOKAZl/xk6DrOmNGWKrTJrjigGZf8ZOg6zpjRnsx8IJPpLDslXIYXjohkw9
WCkk2x3L/Zvq20aKQzSLAkZ279mrbSKYzaSnePRBjulf37yKLrYBALG7lhwNf0XOmUjgDyiNK2gzMMRMS5S7HSJIKl2yHXRj1pYQ5bfGrIH/EpVm2t5pDH+0KaXMLopd
UHIZk/aT4ArOiIJSUGSJmNBUApFsoTZKYRr6p39g7uLKiCbRJr2HgYyrX3ljAm2IH5wwD1M3xQmJ0CgYPmoSqtvfhWccTu8Uy6RbRLYehbgnUVJVGWTX7hWzoZli0iBF
i+/7Sx1D0hFJIh7QwFSXe4vv+0sdQ9IRSSIe0MBUl3sgeDXzR92Fd/6SVRX+Tyrza08zGtfmH3hptm7l2hXSX/UPz/PbpDbwwEJeeJaxDeuaIj3frYsws81ln2baUsNG
ZsDXqra4VlXow6lA/1oPrLqNdP8H2YuQdbQbgxQo9+dzvtNdWKRitceobBXNnTFYgwEyALj7Bh4b92lCZHjkgoUI4Ldufl9jwQ6RblqcKYkafXlRwB+rq7T5T+yk/V2f
49ikr2KDHmwGGOooje69z4YtpmeY7zYwee+WkEkXie2/t/jpRyYiISNHC5LGpRZezBuedGh+rFirRfE1vhxvcQHE7xfIMKKDCpigK7+ZtPABxO8XyDCigwqYoCu/mbTw
ihdatI34yFazXyR2duUyWZQLnqTY8jDou77JEEoB0GNYojP1D2/DHhHjjZNzdsmvFcV2x2jP3h4eQf9uQll5RwrHmd9Nn2eLxq78flu+VUdewitif0xUKqqeXidp+60k
XPOyDk3IC0mk6GbfpWB41J+G45UZKTl63yhqYEDROyIQ5FU7qt/LRBAl/0xMjVt6/ArxS/Z166l2bwIqCG9P+1YMOcUs0MzdPEirj0jsMEvO/mhxDnDvxUZ+Czb+iRwj
CjLxQUI9gizqOHnqSzXOtfYOXjc2w1gU6tZCQaytV0oZKadloSmWDBChbLy7Sskvb/CtFR2CoZuCGD1ddwUCPjFn9ltI1BGH56YmIhbYY2ZWjegH+Kyhta6LCZWrNoIS
f1XmWeKMuMWfg7yuQhFDZHCZH3csa6a9gdALA9kjGgap5xDt0B0gxf21Up3N66HXjB7j/ebJ4P9Qol87BPW3zMqIJtEmvYeBjKtfeWMCbYgXIAyFJEShVYYA7MSXw8FG
OyeUn/V0bi0lznPQpKpsO8qIJtEmvYeBjKtfeWMCbYh57mVJui12ZNdKUOSsQEvGo//0q5ee91lX/axB2xiz1gaLHStM2VqLzUS8eIkL95ydG77qT0pL/25BPXQ9DqBy
nRu+6k9KS/9uQT10PQ6gclOjHu4orL2dyHs7iQpZJMNdMd8wPZHT3ZiEfm+TVOAw0pxHPj22tGigAByBayUfCrPqzge+g22Bp+dJaQJvBsAeUHOXnzq3NB5RqCXbtZ9G
MDunq8MY4DrEMG0z6ci4RmxKVlVH4eDW1Ah1R/vCYO5mu7yWH8wg5Q/j1zGMCnM3AuqaYP9dGDNE5NO2TwaRQCYpJYsN0pmyBFSqKQ78zboeZwTMC0/rBJXC5QKs6vNw
9INhGR5EwmC+DRGHS4zoYCfJ0y9/BFkC/5N14HFjK1JbGXUALXTyia5idSbav9fvoPejuWTbTvma9Hj0YVw56aD3o7lk2075mvR49GFcOekKJfO1cfok5qPGDTTPYnM4
9uPCM1s/WU4M0HvGzaK569v2yrZbIQCHY3y8nboRbUYU4ThECmfSFye2QBoBHK2xgCu5C52dkTk0oIJV3VKhtVzlEg4dyKqUbMF7Ol0dzqf8CvFL9nXrqXZvAioIb0/7
48tMwLZuIDE2TSZaZWh4e7WAk3mtmQzRuMA4kuAotOT/EpVm2t5pDH+0KaXMLopddhVLu7R+F1+hkhxiS3UQ2WXukBiuh+3Mtss7hLjaziT8y7hhx5P2B/5q0km5UAv4
8b0qqSjGDgcV77iDxmUsdPG9Kqkoxg4HFe+4g8ZlLHQ3igkS2KentHmRoXrIcECCLXFZptCUdj4NUXQPRtYlM9ica4RKVKf3HzOQaLmYxYL/ALDxn0rDA2liWlB5d7+/
K9AvsnC6x4Nhv5JNDOdypFIUYS3nwLBiPBfac8ADFpO2QrCgF5QQKfvLhDfLa79xzr0PpUFrGHIEKln0/UyEG6CKbZpJmPCZqSbis6Gv0v0X9Wp1kRFGJC4OA02q53sw
yogm0Sa9h4GMq195YwJtiE/vM+op+bAg2mTe19y28hUANn4dyaPxKREy/F6jf7N51hiKIUG3Fvfg731RcNZO6ewvQDNHWcHejpgffGmvrETKiCbRJr2HgYyrX3ljAm2I
uOzQXclVuvqiA8zThjIP6smyMVRYE3ZLzerOSGfIZanj2KSvYoMebAYY6iiN7r3PElOWUB27D703yAvI2cWR3cwbnnRofqxYq0XxNb4cb3E2hfdp0n4Crqjvl0XxgxMl
TdkmOA362ch80eQ2wvTPYMqIJtEmvYeBjKtfeWMCbYg35uaVbltHE+5B+JTx4SZpCg8caiE//oiZJLTh4cU2Cx5nBMwLT+sElcLlAqzq83Ca54B3V9Kh1uNe7feE5RlO
Wxl1AC108omuYnUm2r/X75x+3gNqZjHtnzFcIl7CVJW7q1BwCVmF18KOp/+9mELGyogm0Sa9h4GMq195YwJtiKyIjzKymWve6oIQZTlfV5pBPJGjXtKWPbanZZ2F0SzX
Q4mOrtHm6PtTUgVFJ2+IxvNV3ehRcDckwS4SVSEYyqbKiCbRJr2HgYyrX3ljAm2IMqQ6kWSEYoputIYJzYd/7Aw3OYwJ2IkPUWKW8E1o8Ejj2KSvYoMebAYY6iiN7r3P
rcUhcD8sTuy83mwg2Mx7RcwbnnRofqxYq0XxNb4cb3E3M8zqhk60ZVIpG71xsq6+sYfZvF8WR4ZNvPNFg8fZIPYOXjc2w1gU6tZCQaytV0oZKadloSmWDBChbLy7Sskv
Rrb52KDHDJkxcvjiiU2eT8BxQBNES/U0OWbKWhwjZAeL7/tLHUPSEUkiHtDAVJd7bLzFyRvUC0wg/SUEbrn4h+Ap8bqzYUiqf18RL3gPuLRCr+NUGaOl0kwSVa/A22O1
7BuwCX2V66t22M8YAcNXI+mDcBfe4IEXlKVoADqncd1/QXQAldk/itQXYx4BVOdVBUzX/o7ivPNL8/I3T6dDcD/PjBJ74yssMfiXAlToDeDwCp9UpKSP1t4y+0eb8lEj
0z/G+h/HDknPxs00mfU8xgVM1/6O4rzzS/PyN0+nQ3BnrvOYhPWjjoIJNFxIK43svMwktjqcHHeZXHh3hmai1s5J/EmzkoiOcWb3CmvI/8BX/Yr4Ly7ww+MbVhLn8Pt5
YY8oo6Tmbvg/IZFVRiilvLzMJLY6nBx3mVx4d4ZmotYUjy4U+VIPs2FDcT2LyXwQBUzX/o7ivPNL8/I3T6dDcCtoRfmFafccscg0n+/OyxWHebJy94gnGJHWe9Oipula
wdJCjvrh7hqmLAG/AGcnzY22yYjwesoun49t7+9VtneVyqqN2PBJahZZs1GzWtNivMwktjqcHHeZXHh3hmai1u3nknmm4OBYOonpNALd676NtsmI8HrKLp+Pbe/vVbZ3
frV3RSkAlb/j0qCUZngnGId5snL3iCcYkdZ706Km6Vr7dJ07VD/jtdjsWxUIdAXhBUzX/o7ivPNL8/I3T6dDcPuh5/+f4hB/AZ5fZ5F6W6PeZNcc6jxwJNX1NA6UMioh
0Di3gqF+sLybZbMGao4u7QVM1/6O4rzzS/PyN0+nQ3B25I95xFbLS5RpOycc86Yj2lYWrWg6R16ZYcl8uBhxsUa+RI+p/MTikYAt/BxFDMUxn4BboK4jKdZD1JeeGPsV
Y4/lcmJD193W4zY01/Rv8T90ccB6aYcMR6CueqqPviX3wXDXWg9K3Kzh4r993bPkBUzX/o7ivPNL8/I3T6dDcHlUIgB8u3VFCXfgpUK791S8ui/k4lqp+l21Hb0r4djt
WoUL5zH1AyptGG2oJmnx0FHULok0ArOizwY141vVA+5hkwfZ3vF+P86/3RvXvCmRT+pYENSLQukftZdMz0REAMJVKVACf3Ii/zBYVSTt5iO8qhKlFqzSOEQS0wquYo2R
iqMrnjEGJuTBTzy5TMeYMU/qWBDUi0LpH7WXTM9ERAB5i842tbjgb1XKsaft/6mZlRTcN0Jzwz0ize/agZabFIWz2VYcif1dyQ3TIARzRL8tAs4dxocDQJETu1P6IB4Q
00ndttirpnAn3FXM4UH+AW9zWpxqwBRNZZjCbPYAeW/BrLZVZLu993Y4hFs0OsTLT+pYENSLQukftZdMz0REAO2c9GwcitZv93R1v8fez2OkQa4Ct/yuS7OSlyOq++G0
B1Yx2XYp+RtqVBASxVrBvE9YKziAbWW1a7gmqZ9YK9cA+JfoYu4KDzjiehdMftrSeDa/LLJjWvyH30n+kcCOvFXIE1TvahGIEstUQFxLyVRPWCs4gG1ltWu4JqmfWCvX
mV9s/ztfyXduB4W/ewzf5B2s1/+wjuENXuFk+ZxdY0+j0yZRRe8vopIrV6nq/gYMT+pYENSLQukftZdMz0READ6mkQfDmLgLjUsTy12+V+V2G3+LSsJ+ohfeweTjoP/C
77Pz/fFVM8cNueuwy4/klE/qWBDUi0LpH7WXTM9ERACZ1TXPvIkAsdK7FRJcOZzZ5t3LmurhUmlyWasCNIxvYQ+hJOC8eqKyeQsM4rcHrQMwx/VUQ50AFR1219X1QbGW
8DvitVnxeQRNnU+xFHLUlObdy5rq4VJpclmrAjSMb2FtVScNVIATxviEG5oponDzT+pYENSLQukftZdMz0REAJOJC+0Cgn3OFRTItaxZTaatleM/lyCCY7NYCEnKLUnD
0TzqGL1Erv27KrROdSPppEeQdWr5CmrQ4Bj9Cb/Gek2KErj6wDaPZ7GSisuA0L9PkV79jA+p1AVIJm/EhLTALxLMRb9bU6BijuciCXNv8bVU+3rdX8WJsXLjZ1y1Zfja
trfXr0S0iPm6dmTRE9m5LqdW27l+RpXb9KfuydrplGj4wKZucswBHhVsEz8CH3ja277X0ZkOxbUcWls/kDYNqvGLxF3AJyF4IFHPHXeCOOwdglqrDLQbqsf/8CsoUl4Z
copNJGEjOiL0lQBr7tGc0RH7t1g/FNoB5dgeqiVHMruLNLVo36CJsO8wQ57oL42+nHGDSaj1hAVGl65Cz2IA1FHFpfXZ4nx7roSfL+VBryPmYZrzgb/FN7VovGbra5Y8
Uk0Xo/iOORytKKgvvK7Rbh2i/wE4d0j+T/V/aSo1cQILuGi7AeipO8Q4p26jTfU0zjMsJqH0M7jOWK0cQhQNtkfHIoxe9XquSEvf5t0FyXwzzIlOZVqo9kKAmco15qLo
9Rcc220qLBp4zlPu0RRUXy+GRhulbLqHu4Ho904vjDqccYNJqPWEBUaXrkLPYgDUdJnYVqV+LKtbmShesURnbG2ggoMsjkBwPrhRP9KkgGfIVeqrava89a5RAPzd96Sf
GhKppxCJDuHAaLblceiwDKfMD/1iKQzzgjYqWLg3zq28gCZW2ghDXdsYo4PGkYs6UdIv4pdEiBf8L4nokRjwvsdF9sI/soc3XZSiL8Wy2XVhkwfZ3vF+P86/3RvXvCmR
SW9NF6CKBuHLdrfZ8dEq9nUX0M0Huz1n/2FahbgtrOcpLIB2sViVJhhrYT4vIhsWggLOmCPkFgXqsyNh1JZ0hWRCrLYr1iNl4IfUMQ/Yqv7BhxwGOXvFTJyKCq1au/3u
DlnCS4SR+JHwqj0zdMRHHWRCrLYr1iNl4IfUMQ/Yqv7uUEzQf4UU7gvhEhUjK+KddvGYQxlf5/zvSRrjJpslU0lvTRegigbhy3a32fHRKvbD2Ug3sLNMeSvyr9au4PjV
7LWYvf12qIcwIVsTnQxdFAicC98iNqFyFhP7zaL+Qbc3PxnIhG4enjXApC/sLJzbI4/wSoU2uO8GIVJC7em7HevJBKP6AZtMHMHYlkijlIWuLO+vk5M9FpJrEpM5cq/x
KawvAeCWDMk756Lj9NUxEGLw8EONRTiCKVwTP1lZJpWuLO+vk5M9FpJrEpM5cq/xDBhQnGZPjF9XchlIjvP8CWNtKVU6+ogXgNc9s8+jusZJb00XoIoG4ct2t9nx0Sr2
ftOVhLEGDXPJL/nrqvEu+U74YxNnVR8aOqIx6rMYdJE4xfmj4SZ3Id/joEPVC6HoJnb+7shUuLXR521sn6VFl2RcNwQ7ub5FuxILF2M1GMq/RVcMyqT+aeKzfmzaDeYC
kszkR9DAT8dXxEBjIyTux1Uh59ERS610z74PKFcPQirbhz7dQNpnag0SBmEdCDMeu+Xuw/Vm7dEqp+ZVh0fU6sj+T5P8di6XieeA1YJl3frWjw+XAyK0VB0/bjMAmj0/
DAReEdF47j6v1kDyjg+eBp1gOoyi4GCLsUE5eTueqihTpuA7aHOlUzvSIMDFGxtbPZQeFE/k64BS5TP0mELmwMvCUc90x1uyyIqzT3Pxc1aFGq6J7zMN2VnQ9q9tZXSO
RK6q0VoLiyzL4hM5mmYYxwnyKaneo3NdPxy6khV1/A/LpK3sKcSvezoVff5r3+M1e3fr/wHHUN7KUUH5ZmmYLuciDPTnZZazCr2nLu1ibwvjS3BifyzZcRp7QOKB2kcx
OphwATLtaA5C0EoIoK1V9AHuVfRGB/+kXLeu38IVCAjnIgz052WWswq9py7tYm8L40twYn8s2XEae0DigdpHMXEHFErppmd2Lz2lv+fbEYhisn/Lycxb5unrp4oyTD9k
SW9NF6CKBuHLdrfZ8dEq9qQgLfaVW9wip5l5kSqsCglAt9w3BZXKqVM8UkrHqlw5fM1BrTDvqCSawc7CNQIQ/0SuqtFaC4ssy+ITOZpmGMcJ8imp3qNzXT8cupIVdfwP
vIAmVtoIQ13bGKODxpGLOrfR2gm4Zl6IrFrrWt67doUCH83vxX/QWNq//2crN0inMoZWkBLm7hLM9gRwhbEHw6Gndyn+oG/l0NLoTzNfO291Ft0Ka2eY/nnARyCrL/I8
PFBEzn9gg5VAfcaQbcTD71s4KZ2JkgZadewsAybRpfvwnLEC3y6LNJ9iQxtO8tTJZXl5NE7y3esENohEMAvcKtOI/BdsHCMYSJCpQYiEyLA0s6/XOidH1WbxPjqpTW+h
dxu7Zjggox0rnB+OyXID9tZOsbEkD5jHOWvo2lLMEFJto56twzD80DlDOM/0+xuiQ6pzMPWmXzK4zGnbHWmrWSAVpob4eDr7T9xB3v2u+jLYfQxJpn/EsFoIdGQdPoCw
34zOlSU+0X7tI7LXb0XLLjOw6DGRUH+IzLnjhFqhh3+H+Qr8TcUehGvK09xqj+SHlinxHmI7H7/VzkpfTqR69Opt5fYFgXGhC/j93uCfMHHBDs1rcPBhsrx2FFHTwBJQ
h/kK/E3FHoRrytPcao/kh5Yp8R5iOx+/1c5KX06kevR0azKsEbD+cRFf9WUBP6uNZKP/2CPuEaVD6HT6CRNtZVmS2/MevkzUvChwixCYPsAVKKapEo5djxxA7ah9S0VP
8uYii+eA6wh6vGPl0c75rp0hog6ZQERQFY6yc9IV7uiH+Qr8TcUehGvK09xqj+SHlinxHmI7H7/VzkpfTqR69DVkTJrLzq6VEDuUEtARovSmW6vIoVqss2d0zovJGcst
/YgiSz/i/Eu267YIlzljoMmHtMaA+RilsMAeNqM4HYY/n+j3daE1BEIWnlhQNM+vUcWl9dnifHuuhJ8v5UGvI2Sj/9gj7hGlQ+h0+gkTbWVZktvzHr5M1LwocIsQmD7A
FSimqRKOXY8cQO2ofUtFTzqYcAEy7WgOQtBKCKCtVfQB7lX0Rgf/pFy3rt/CFQgIxhcW9VkrD8zvdb6W2qMDbhO2t/zi18LzlXuyp0bXINayLOShbffveNuG0SkkslFv
MWEdcriHeqoqXgBsOX7XsTOw6DGRUH+IzLnjhFqhh3+H+Qr8TcUehGvK09xqj+SHlinxHmI7H7/VzkpfTqR69LLhoGOLpatml9mCgyzNYSMniTVigccbewb+BB9gt5kJ
3407OnK/m7nvmPLa25N2C4vUqGZWqxajzZDkGkapTK7x7Y3XIsE7ImoF9NaNBynZkm10U8ol1VXeEYkGLXn97UVFaeHXAP2NH3aA2eQ6evbeR9lZuxv6P1FYSic54lDb
fWi+N0fVx4uytpEVUHCvp7B0+FN6qoNgsUv3h5yZQhhuWZYEpfHbap2Fsi7ea3CrDlMNYa5M0aXxpvmazRhdgk2qkMdYaSMzvzGgzrttqa6jrGurm06RmdBj72gdwpUB
I7CAHylzkk3ZvVV34r+i6a0fj5vbmf3YGa4kuG/UP/qUkz2mEv6oiPkIrn3uo/4DFjPmkFFofbM0PCXpX1hekLBLzmsin0b28WoJl1jInNOhZltutuyR8TYjAfPduqo/
GsQELABHke6Xmz+4TMbRIbh2xNbB/9Xo3/bgtUcWlgvyn9V1FfbwNpIQ4T5o9kfjfaFDGz/8ymX35rye4zfE8WfF2A1gpy6tIugCDgN0ssJvyI/9WwWfJRzS3Jb8qoAD
9jQetlSQy17R4CYRoN+kRxRNp90MIImCrFgEZ6I3LKiBDEiH/InGj0+vk+gk1+4/SEORe+wb1w2KzqHh9M7CB5GKp9IhRvF6A+KVxeQWfPgHAhf695+X8e4QitOGqeXf
Nb2rC8dNjwqOq3VQWYrrRbIyicF9RseNA4fwLZvfTWVhmbRyOBTh9FztLMINMxEpNNOGVzSYogROy0NuM4FnBM1usnL/WGf5ZaT99OcUppiLtEp2RZrQ1lOkdvSonD2Y
b70MB9+3uHr0pbrY9fkGnKp97GK0O9QmPcjuL8Fsiul4IzZMAwgy6IZvX4pY4RWn0QDctXE+W9jxpRNlBPzqzbwoLoSj8Ch3KcYC9y2UR2HJC5EH6oS9fM4/DVgc/nPA
poeGgE3TWSqHzRSaUkGSkW3kj5IuwmN3h5DLkGKb/BVrqHxya8qOIiv364e9br9U5yBClhG4PliWU/t4d2tGFaY4FaJYqKM/QU4pjO+VtA9iXwSqpNOfH4lj8DuGxmQQ
rIuexBUL6rcz52VTxo1s+BW33nLjYUPFXYMrIDTcmvO1wz763vulT3mf0ItXqIltxiqdcNQeFJfbQI5pO5FX7CPREhjDnZ2NjZgxKrboNTja0ugNoXWTULyaQa0ogQ7W
yijZh8LmwfiKibX/WkCyZJzidqvHNiqpzuaRkIh3gxpkx/BKJOOGTBa/SaAH4ckJZiPOhWuHj82avCQHacBylG5p/fmGqi5f9yuET/1k5KkpGfi0CFcNAq4al/cucQ29
Yl8EqqTTnx+JY/A7hsZkEKqaDIEn01S4utfqdfhWOLwRx5XWsaZ1P5Ib+cgBQKHLzioiWg16mApuqj3kgOdwUndUlHJ2klnYko+ZbKQ6GJ5G8bZGCqjece/g/FivvUmd
gq+KeA3zsQFVJssfuOiLMJXKqo3Y8ElqFlmzUbNa02LCjLpvSm2BR20EoQoq/teJfNHqd942fE2Kycf84VudnM7hHswS7ovAuBePsbrL5+1uaf35hqouX/crhE/9ZOSp
1yF04dT9+n5mrGDngPjxBFKQICoT5NXh9OeysFF7krhuaf35hqouX/crhE/9ZOSp+3SdO1Q/47XY7FsVCHQF4Q1t4q8u+fJk5s/Hl+9AWojSS9H/nlBrfKw94zJIL8wP
4XUFs/+M8KggGJ72bQFkxM4qIloNepgKbqo95IDncFIjawvji9JKH0JvVcVZQXg4PFBEzn9gg5VAfcaQbcTD77UTHCpSQ2aslrerW2UDZCY0itBjyCorvTWpGUW70622
DjjRLCtJYeabQ4yDcoJQ+USA9qTPGHOo1Z0XW0DYeaspOsKjCzPm1ewlFzbQjbrl+e7PK+cRFCrP98CZvANUNN5b6tDFtNM/4Gd9G2x59cpxxiZ61wVbcxqfDgOym4Pw
LVkmdhHzezXl3gwVboahydEAe40MOUxvivZFnliY92fOKiJaDXqYCm6qPeSA53BSYiyQv03aWLDgCet9vB9bxGXVNNGo6V6qC03r9zuxeDLUJy66FSKqpKkQn5j2fqnS
mjW/OCp7rpilyiQ1LZ3o0kbxtkYKqN5x7+D8WK+9SZ2Cr4p4DfOxAVUmyx+46IswfBpnd/B014ESoaLSsMz5IiPREhjDnZ2NjZgxKrboNTg/fgpgL3gjq5BovzQWUWgI
q6CiEV2iV2uMSQbYjvWfMy+ha+klNnElFHPmu2DCw13li6Wwm7GWWpkafS/qwSADSjG9KVkIzIbAn7+A27qNu9d+FmzdnozwrEFseokVkY8319Md2NXH/tm/NIOPmXGu
ITvOaUXpn5wp/GySvq+pzDUbphO6vKXQT6t/KCilIcAuagRZxg2EwmbPNyqM2OhWpS3CJ/l7To0zyoloZbzI0uU8bomCKLqu1IVVPRUfahVQHiH3V/jdPPkwE4KO4qnV
8KCxok2gA5OJVZrTd3rDTWa2aeLlJv+H9lv7OMaCDmyu7bi1rt0o4fckyoBexE6CWLH10c+oNwXVdOyK+S4EOEVFaeHXAP2NH3aA2eQ6evZ9OwemgAmCXpW+v56s3ysj
oIg3PiLJd+q/jU3e2UJ1FySRZ3A3MHMDQO3FXgmmEs+BlE6BxAFWPglDFf0XlEDYQao8ZV5M4uh6jHiP70pZAWTH8Eok44ZMFr9JoAfhyQlWDwOm/StrULS6Igm1hH6Z
hKVEqQB3j9JqwN79R732uL+nGLOmT8PRkhdc/ba1PhPpBZDnOpaTc4WdvrzZe1cMcOjNyxwT6PAe9JhMgD85kVZXw7BKBx//sjO6afZMjXXtyNwyoRM+wLZ3Y9mI/Qvm
d3ob52tYMj2hEDvRAptNHyZfcYdpuS04g57jACPfRzBhkwfZ3vF+P86/3RvXvCmR/YgiSz/i/Eu267YIlzljoMmHtMaA+RilsMAeNqM4HYY/n+j3daE1BEIWnlhQNM+v
9Zykw6Rn0UyyqVWyGNHfls7hHswS7ovAuBePsbrL5+1YGZyUowpZpFCWhtplQ6fcw24CNW2Kf3yAc/afDNoctKBtcAjkJk+lQ5nMC4V5m2Fyn0EB7W1neic2RU7pUpJb
PJiSp/TammOmvl3YmqixudQnLroVIqqkqRCfmPZ+qdIxV4xc+kN5rsyFpTZOGjHNiFvzHtjCimZvCUI31lkp8Bo2pHgdGSj26xvjyYaUSWOdilUfYvrjOPFix1CFrISa
eXrLOFUuVxe3GKiGQHSH86Vwcc94E+fAqbImtGqOjUAH5Pvj5669mfbRer0mHKr4eXrLOFUuVxe3GKiGQHSH82l3ClOUs9B8O5WngBNEpC1Q+15j50kSN1dCbZ46oTyA
LVkmdhHzezXl3gwVboahySg+vrW9xFhmrvHetGFVZI4dCcthSW1nVe5P4Z7CgX0TyijZh8LmwfiKibX/WkCyZJzidqvHNiqpzuaRkIh3gxpkx/BKJOOGTBa/SaAH4ckJ
eL6gdpi58j51v+FOloxjkVhI7gkMXnaiGrOjJFr/9tVyn0EB7W1neic2RU7pUpJbPJiSp/TammOmvl3YmqixuZO+lCBL7wwwTR+vMtdngtkffoF+YxsPZMRdl3TP6Fgp
4z4TyBvythcHb/wQDGr53qmtAxvBqmFlO0ATy8GPLY40cufLfMklhJWdWfegViXoirvrfLG2AAxrmt3sx757PQ7LeqxQngvS/C8AKs9v3t/GFxb1WSsPzO91vpbaowNu
E7a3/OLXwvOVe7KnRtcg1rIs5KFt9+9424bRKSSyUW+hzjSkNsNYQwWGRDl/ALjZy+/KBcRvy6e+qn/l5K8lCvAUubkiQyO9B3/cBfUJmOqPW+wpuBD+vbfDYFomlT1U
UWAjewyqcM3W3qRQRNF2CqRTog2q02BB5qz+r0mHagtibuDieN6/6YLGJ2h3d8ySnC4cMrskBoOJxz3lFWu/NUWFrcGo78rqdTk56/PGgFA40Gg2NzW9lL+w8iVbMl7I
m9GB7kVeOqBh6Ki6arh0WwkFg6JflAEtBx3cj2sWsQ7KoDXDvRjl89SXhun75Fez/YgiSz/i/Eu267YIlzljoMmHtMaA+RilsMAeNqM4HYYOefVOviyIfJ895RjjlXDI
s+rOB76DbYGn50lpAm8GwJmpK+M3fgCleFvDwqL5ED2H+Qr8TcUehGvK09xqj+SHlinxHmI7H7/VzkpfTqR69MukrewpxK97OhV9/mvf4zVc87IOTcgLSaToZt+lYHjU
tCFPb/+p8ZzQoDpJR9Ie8dA7Dinzv4UkwnEUOh5C7zqDRnlTVCm/lSpagxjWTRu6Sovp5v1Q/Ic8eGjSVSHx5F688IZ2/yDx4uryrQ1gfyRYGZyUowpZpFCWhtplQ6fc
w24CNW2Kf3yAc/afDNoctBEyMmh5BjMlLRrMfgNF+Z9Hg7h+EAMrj85zck+SKps8j9KxeZCHTDtVrlW+O96HOHdnZOt2+LSE0GzbwZ1EoHFUl/x8w85q5IFlbWmOV/FA
m+qjK8OCr5cnlGLxzodoXZoGCa5kSQBKDk7N9B5yBeb57s8r5xEUKs/3wJm8A1Q0jHWGwBtxudoCIJMswYnSvTL39MVAAOyvgV0+LoSE/iyNpXM0O9HsYEpA27rm50+W
B5Go9LH3StQUC0XBYwXg4C8FMAY0F3ES6XLEY7WVfBI/r0PfKUnsXxx/HniBsHtZ4RV5gG0ei3t5gVs7eUGIARW33nLjYUPFXYMrIDTcmvPL8+k7ItaYXpDgPBzZNm/N
90Ur50YUlBE0Eozlo1P1hHSQC5vfaCZW1iFACuwqc5iww9DhfVo67vZkJX8k33V78RVBKHjHqRUa/h4+e8xRyMODxBzBaUj0w2z5q5mJ2MQm1Nc+cdEUcbI95d/B6v/b
DXTI/qFyk6HD2M5GyQHoJwU7tcd8JUvmpWY6YwI4nrHN2zbtICS7LPpyY3GIS8JXxohr1QGDw4z65pOgg/RmARYz5pBRaH2zNDwl6V9YXpCUcBghtX6N5mWKF9glTrXz
pC2WC+rken9jA5fw0Tn6eXQwIGJQW8fNEM4vYseNPF3b9sq2WyEAh2N8vJ26EW1GW1o2mawwQz2JEVOIm4AZB6Qtlgvq5Hp/YwOX8NE5+nlGBih6ma4OzP6wshxeRiVk
XPOyDk3IC0mk6GbfpWB41FqJXwrppvicfRiEIzHdmKO3mLTKbcc0HE9Vu9+9S4KqBoU0VLWpCgr+22kEgXxmSOEVeYBtHot7eYFbO3lBiAEBWNpsrXDElIcZHXhKFD46
pIZdTIdkv4A225Sl/0sY850bvupPSkv/bkE9dD0OoHLWtTuQsY1F7+wJCfO9Ql1h2/bKtlshAIdjfLyduhFtRmJfBKqk058fiWPwO4bGZBCqmgyBJ9NUuLrX6nX4Vji8
4AioOALzHftNrlkokhs212JfBKqk058fiWPwO4bGZBA87l5H3MgNjMIi6n/VH8EFmgYJrmRJAEoOTs30HnIF5vnuzyvnERQqz/fAmbwDVDTeW+rQxbTTP+BnfRtsefXK
4JqnN+kfOdBQc42WY5FktM4qIloNepgKbqo95IDncFID/ioxVKYlmwMh3+PyNfT1FkuIuzbFohy7owv/9ddN2Fzzsg5NyAtJpOhm36VgeNRrqHxya8qOIiv364e9br9U
5yBClhG4PliWU/t4d2tGFUhaBR3YW7gSSlA7v0WX9uXjlXgRAl5O1VcE7KFwenPUtRMcKlJDZqyWt6tbZQNkJutinWAb4JQk7Jb+LASruS3R5ShRIl94UvBsC1M5FJnJ
VbVFLK3ISQ+/Jb0VFly0LpJMpxiOh+8fKvqp/YZ20Sc2Xtr6Wpk9OZJaPXEOX4MWVbVFLK3ISQ+/Jb0VFly0LsoYjmxmyd1la4chz2HdSolMNmZBj28HaG6lRkEA1F0O
5Tgu/xB6F7GLn7KVYhepQi1Tdo4pgIva8/el8GqzUHlBd3zuCKbj0ZGQX+Q64sNVVbs073fcvrxbHlVKp5CWr17B6WZSmR0mtH73MuNXfjlLQNa/FhOqWiRREx88UrqY
lM9LFDk5XemfePQjdp0FiCyO42Kb3jtfCEhJXIAZkj8vN/QlWkVSpKSXXyM/ACXJqa0DG8GqYWU7QBPLwY8tjopNLtJRAGAzZgdkVxQc+Wp8QWkkz5pD+aYCYVar2C62
md38PGjHZ8sclBzaxAo81mcWPM93BzVP44jjI4xjzZSWy8KLriGQ0G+4n989eBY+PVshldargUIN4vBEeJ41r/wcHRaRFkau1L2pP2HVWnP8CvFL9nXrqXZvAioIb0/7
DCiRfIsqa7ChJXfuOvabIJA1vXO/qJIf+eZTvUj1RMYP/nIFXLtJv763lmQ0t2skMn9srzx+7NtMSagtmFerbt4PzRtOedxQe0z3JDxrLx0sBuyk3kLeijTKUuhQgG3j
09olWcmo6KxTyx7ZpjlIthb3duhF0O3P2gcOryNh0H/gFdd98i1+l6eWkLsbMptoe8w9Q6UyQgNAxQ+i8Bzn3eGZMSz69250nP6vU2tNa+KO7Qp8yBHtObE5CTEtEvkJ
ju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJju0KfMgR7TmxOQkxLRL5CSt5puGT5o6cnc/MlCCVU2WO7Qp8yBHtObE5CTEtEvkJ
ju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QlQDpc2VOLGFqGgM+J4vNKy
ju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QnGwSngAvzjFvW7ArPwPXyc
ju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJ
HIJBbOaM/2WyW5EAIvBEWY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJ
C3LXETpH5vPlj+YJ8MQ+z47tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJju0KfMgR7TmxOQkxLRL5CY7tCnzIEe05sTkJMS0S+QmO7Qp8yBHtObE5CTEtEvkJ
ju0KfMgR7TmxOQkxLRL5CV/XLp02rKGl5LTwDMFj40zYGwT6Ye40keMrayrlpAKeyu+0QeiBLalTkNhDQR7Lcfj0m/ZMIBbRhKP/JcYafRUKa5u4fv/3HyNCHWUmPxVi
Epm+eUBzFsZO+W3gBFjYbY5IEGpaVZsiZdTdUyBDFXxkjb7owkbC60XvVJHOWzyUmv7VepMByIX73lGdbu/1ib3ZfzNe+37SxUQSZfyuMd18hz4sViIAFjhlAXnPznmY
sMk8sN2oIOWj79U7zz2eZ/ifYfiqLxgTAmEGvzI+TvcoDToqAkJTEKpA/oBn7wJbQi1mAx6+NF8/O4ldWjrupIJXpGJrU1ZY+t6574RPaS1IFGZ3O4WkvReJmz7U2PBF
ov7ywEBicN5gAXl0VWOyEn7Nh194QFWZ15+NFmvR7M9s1PJCF1naFak7R35td5gPfIc+LFYiABY4ZQF5z855mCtA64Sk83XxGDNpApDpjZBQ4UnBkDIrATBm7se0jqV8
o3RwL11tQ6uNoUScwbJCZfL1tJwQiwOaNpCeX+JhXZgbZl63PsTN2dD5cTkfeYM37c5EiR43am/aPWZ6c/XZBxCJLOS+HkbD+vejgUAUYcEjqFdNS+/ooGsJ25OPs02G
4JqovFaNj8aKrBxtVHXv4WSNvujCRsLrRe9Ukc5bPJSZDzJN5eu8D08jzfZreAofyLVZQN/7EUHvj2i78gkCc1zu4R55P3bgtmlTrXX1nobSvTjLV9nanYcA/TEMsmWO
UOFJwZAyKwEwZu7HtI6lfPk9sPRENrFm7v5eTOEuegQK05Dj4ofqDwb4GzYDl25vYKy92zq41CfdXIHHgY0Ii47buKpHLWqg0p21Qc1R2L0H39EmOMVMnxKb/oAbdJxx
iydldj7wohBhDviqq1KbUPQJwODzHsfOtjlqSUfR/jcQiSzkvh5Gw/r3o4FAFGHB5jPuEEYOfNQ0MOenH1KTXQhQXfp0KjX5shmCPQhwVOCAUqHQTa7h21GH6ln5Ld7e
sJqzDo8wrqNbLqJzVPwfPC2hic73UVO9r+HNVhQVpaeQl7R1G73J1Kx0A556GbKOqYNUEi8VKCEejkUbw1BZY/ifYfiqLxgTAmEGvzI+TvcBTxFJapaF8alBcKHqnUk4
9pSOuY6V7j/LoSHl4plZzh0PO8KM1PvuLY2mOQA86bx2DaA4TR0/84pkbAqyspAyEIks5L4eRsP696OBQBRhwQx2kKBOqdgyqGKhGKOdf04PUosJGprncSl4lQ5wpG5G
K3LAg/8tfQCC2K7s7gi0Jxq+mU2iGErQ/l1x8Vwr1XBQT1Xing8QDWY9o+qp2xEGfIc+LFYiABY4ZQF5z855mNfWh+3HjwKujGWwvEkUAxAfNr4vDgRR7T3EYgTjq1rA
t7gCxVKMx3wjGfhcJ7I4sm+qXaXBsOHz5sXSM3VIljaRm/142H9RJEZ5+BTtlmRapLNX0f8rUrVM8Lb+l2BtKLok2V2dIruPQbHyyrffXk/Nzqr26LBZADP7KUNUK0Wy
UI2s516oWm+JWkQsHu7MuXSbgQQb2ZUnXt1YTk4A5n/vSjTLEQ0VHYghnqgK5wEk7Izs3t1UIzBjFylBD1DzKmuOQEBPgr0W7RC39cz56aLRXSmZ5Vja/d9FBNZ6K4mH
6YSRWej+XfI+7Mb633r81uEn8a2nOmEQQUvLv/ScFn3DQw0SMcapIh+7L8fdiFCQpXKHsJV0YqrkbXM/od8iOo+ek8nOq2patvS/rsdCRTG6JwSJ2FAyi61lGdA89DaL
nmFo83c8IazQxWNbcd6dvLqLtX5nTpqFgdPujIvjJEn/yvZHmNrFx/qj/WS/qT/5tVlxfuXrIWuEIg/Q7cCswj33UPW0DBTDew0oJ/lVhnKolGVKtK/6ceVvqkGCMmBV
M96cgFrEe1GbWt+J4pd/RS2jrh9MKRR/MCCJBwfmDpuLJ2V2PvCiEGEO+KqrUptQIJKf/MM4UrfVeAGYMev0wA2gsUZ+ctqxBxL/aTMmaosYACG4zY2L2h/IN9NrIY8u
rXkybrxE8HzbQuWPQshK/ZUl2fJT8Ot7wRMN2b+G/5sSR0DbbdV14k/No9x4SHjFE9+4BAOMlIlNuG1q3DJWkFo5atVqlH38iDZayGtY00olILWknr7uhvhS3wFmV9Sb
hb7NBUMJAj5WnkvUVcUuPZoKXAMBAKSkmI5XHSZdukqn3KQiCwQtkh3XOKqAK0UvLmKRiI2lIu7X97POMWrj67PFIl8/EW2vLIT/kPBcIJJN6ziUEYK9+ZDkBbwd361P
WTO0+iInBHI6QRDVSWUB2oMediYj9kbY/vgz2q/QSHqwv6XmLGaU/dbkr6ra9uJnamklj63cDjm3BE6JR28RwuLOuo7WG0IphdqALh9mY518hz4sViIAFjhlAXnPznmY
xR5+20k+d1ZffvLsAY93UZvYE2HnlNCT5vyDAgXs0WkcTq3V1MatJieCvrOwe9mLMXBnV1+VP+JBrAe3VPQ+OzkJ/s9u7Gk7H+f7wRicrMbqlT/zqrWww1tazcy37rjy
QefJz80JEcPcQP4gPGU2Kd2frUoTqVGuLRCppXr8f7zuFaOw5ZwxNbJo2jj4tJb0ADzOLRIyu4mLDebjC4CN/CwnF+mw8U55Qwi+nPaaaMozlvkAc4fkfgjxuWOeVCj0
HQ87wozU++4tjaY5ADzpvGkuq02dJxnAA0bBUeT5II5YuTMXJxNehD5ZFVloIi1hGs1h8RIf8KJ/apg97GUBdQy+/CHU/ml9OeSkVBCHNc9j4psmSUfxfVvaN6ZTTV+R
rUGfXaxStsferh2N+4yt2mo7zGXDgKHP5rlkvMdzIWlc7uEeeT924LZpU6119Z6GI8I7B/Wnc6T0TKqQC76rH1gF9GkqvI3T532KH4N1qB0jqFdNS+/ooGsJ25OPs02G
6ZWLfuTbJEdK8b6wMHn7D36YZkr2qoKL/GiQfrEN1/2D/LRwCN+m98OGxdtz4K6iAZJsL3VUrvxbexRnQg+wjYJXpGJrU1ZY+t6574RPaS2gJYo4/qKdyPuTwzGZnC9v
yu+0QeiBLalTkNhDQR7LcW/xr2FzC7ioF9D9OU61njnD18hpaarx2lzNs4fu9dsga45AQE+CvRbtELf1zPnpon9nLPqZUkh5lE+cOLxgoHhKwcAM3CLDQFtnnbEt0G2e
j/82Q+n4838fKjtB9tI5yxvO1vU4p9VWNGggz2j83GnEmBPSk0KCZ5KTVBLjAZeBeOrlEqKdGKAqDcSRP2GkN6SRMWV8VsqHZJwFF+bkWR8dDzvCjNT77i2NpjkAPOm8
ntGQJAWtwLT5K/BDK9qURt+qX1+C3d/yg0Ua/uxO/LmQl7R1G73J1Kx0A556GbKOJzLocA2zlF1+59dU0OarwG9nPxYcIBZu+nGsqy4SQD/7vX40qPfgSeaLYFBLjxTi
WiyUYlvx5uAeBWovvljKWwYdTyCH4mR1vvygUtKipZmvXcbxTl6I66xEYpYqkKGrm9gTYeeU0JPm/IMCBezRafk9sPRENrFm7v5eTOEuegSYomhMSFDWD5EQxRsGVssj
Oz4VyjAcg9Zlj+cwFwFDXn088vDiFV6M5iacxke0SJJe8Sb875l3T/xTPlAf6LYcOFsWwgIT/FTLaFuWsTBnfMEuN4kKWQL2jqzj4EQqVtlQ4UnBkDIrATBm7se0jqV8
GJCKhVWPqWAsY4KpVwW9qAyBfM8XJ+Zx2t4lkzABUVZrjkBAT4K9Fu0Qt/XM+emi63xf+m5D8wBOkDxo/PnZtfD8K6eL5NLbMMpVc+XQsMbNzqr26LBZADP7KUNUK0Wy
x9la1CokMsVEgqtdimk+1WTnw29GDmZcozuLu5lWZzZ80/mGpsVujfbjZUh5SZjlTWnZIECJS8dUmztw7jEOTDDvFbO3+L6gpZDZ5IjvnS+C/X3DVnk8QOLIcnhDU81v
WAX0aSq8jdPnfYofg3WoHQx2kKBOqdgyqGKhGKOdf05x+nRKJoZBBpZHiPfBPWW62RSRGFSm7XHFhiZdlmAk7TgMT/ZgCOyrCShkwm8rF71L9I3hoMDbfubDOLS7H5/L
JalJOJpELimcKU9Dkv+3863QmYGIVamwMEu8AzszY6oQiSzkvh5Gw/r3o4FAFGHBEiR2gDb0d/y4CjT7PTh/ikv3OmvGiHh3nJFQ3z/3GL6VJdnyU/Dre8ETDdm/hv+b
ATv/rNjhtPhdYXw4+l0QLL2aZAL08WnD7LMQE5s2xByLJ2V2PvCiEGEO+KqrUptQLkqvMfjvQGi+GArC6JKjyN73PWqsTBnhaWhDWcrifYCtjeEfacfJ8vaCAo1VZBNf
9Fv8SBW1hNzhTF+/SymJKikINysCNi2aVp7J9/SQ+vzPyXAvP+Vj7Z46x1NuMZXVz1hYidLgLlLMRodU25gJIuEn8a2nOmEQQUvLv/ScFn0dpv3bHnuDUaluxzI3Ek9w
ZI2+6MJGwutF71SRzls8lN5SGCzuB7hJgEXnY9u8L3YjEh/TrsZ94TgqG4UqxafvlUl5CRjED9Ck+vXAt6dbtDiM3myTTIanu8Omv/wPmHYfNr4vDgRR7T3EYgTjq1rA
MiMvU5T8ts7YHaviRNyHV2xawJsdGnD4DkXlGP4GTL85Cf7PbuxpOx/n+8EYnKzGEMfNR3w/wVodYgqWdY9wdvmfEII0WDqAqMII/3bTXMh8hz4sViIAFjhlAXnPznmY
fC4yTHSu+z1brtLKeQQnIU+mf2XkDDhoLnYUixGk1goYACG4zY2L2h/IN9NrIY8uUjy0HmwUdcDcRfBV+xnwmNXiwuib4bbcu1iX0TMT/mSWTS2ttOzlxDpWPOxrs38q
ijdlabzK4MRgIN0035r7BVo5atVqlH38iDZayGtY00rQQi0bRcA6cuEtpx0vzzy7+J9h+KovGBMCYQa/Mj5O9xwosgDZjVA0Rp0BWmzY/hBQYv3ueXz+sRW7OCvQ9xDl
BAUNE/A+3DM33955U7wY56Mxc5hCEQMMhxCO7vc5kvEWaHVIKsamXFkZ4iOizUon0gu+0siZgpup1A2MoJfBZeQ9YAZZZQdkuZsFhVVhD3Rk58NvRg5mXKM7i7uZVmc2
Ppf6qKl0W+5AF6mnuenPR2HwPaa8qPI/bWBB8Yt8PtRrjkBAT4K9Fu0Qt/XM+emimdF/cGZeZ6e7nWzViNhy21ObH6yLLgULvr2D9+ptfVCLJ2V2PvCiEGEO+KqrUptQ
jhlmFDrt02zhC++A5Zv96MSYE9KTQoJnkpNUEuMBl4Fv8a9hcwu4qBfQ/TlOtZ45aKgn0qg5MDAxSbjZA8/BxWCsvds6uNQn3VyBx4GNCIs/Aws2qcupguH7bnbpw1G+
UE9V4p4PEA1mPaPqqdsRBnyHPixWIgAWOGUBec/OeZgQ6XS2+NmR7m+MCBi8xWEo/8r2R5jaxcf6o/1kv6k/+bVZcX7l6yFrhCIP0O3ArMKzr2XGzKvKlB0UC5c5aOWk
sL+l5ixmlP3W5K+q2vbiZxCNePsy8lLUARtoAvtWnZRqO8xlw4Chz+a5ZLzHcyFpXO7hHnk/duC2aVOtdfWehjVXGmqBQbeqI64usYALu/Dfql9fgt3f8oNFGv7sTvy5
kJe0dRu9ydSsdAOeehmyjvTszT/eQosMu2fJHiVqM5Rk58NvRg5mXKM7i7uZVmc2LFnbSvTMqaxlpNYM/CWlx/Rb/EgVtYTc4Uxfv0spiSopCDcrAjYtmlaeyff0kPr8
tllR1I8Q9pgmAW6QdM7Q/oo3ZWm8yuDEYCDdNN+a+wVaOWrVapR9/Ig2WshrWNNK3w+NVzA3rz01mG4KfxrWxXSbgQQb2ZUnXt1YTk4A5n+fcMotRVl3VGlpyX7bXvz8
cT8+5yFKN+x3DKItk2FiE1Is5EWTTRCYHHXJay7yL5HS4Jz0K8061v6puBm7KQ23N0GPmWalwTnjW8krYPt0UznupGqaHE11+ctL5I17EHJNndcOoo+PdtvzB61kpap/
T6Z/ZeQMOGgudhSLEaTWChgAIbjNjYvaH8g302shjy7nr6zxeKiIkUFMx2WoIPbP2RSRGFSm7XHFhiZdlmAk7XHv1YRdPEuC7iGCzzfDbXLItVlA3/sRQe+PaLvyCQJz
XO7hHnk/duC2aVOtdfWehrwzU/VUS20EFWPmFaBqX9UQiSzkvh5Gw/r3o4FAFGHBDHaQoE6p2DKoYqEYo51/TjLJDYngC9iSWSp2Y5cAEHilcoewlXRiquRtcz+h3yI6
0uCc9CvNOtb+qbgZuykNt6fcpCILBC2SHdc4qoArRS8uYpGIjaUi7tf3s84xauPryRRsSCFynAnzIKUQJ55CxY4kUWkmnECymLfLPa3Q55TJ2yL9tPwxHYQdi0jpq3Z0
1iRbfwI+9T1KqWhuV2gQ9C5ikYiNpSLu1/ezzjFq4+t4MoPh6dm90XZX1jegsSbJNtXnXeVzf94QRinks/40EYxEsXeVUduvQ/EfAFUla3j5ddCSBTIo08r9EQ6D3+L/
GIq6IS8YdaSN/NhNq8/dvJKEUQ+6bk1aOkKCpoOqwAHCKpDsd9Xff1KXyKTQZd4iC+XgJG957d9t+SIQYSTLwq2WPl3UpB+JWOqJkkljU1elrkfIwh6OxTF0L90GrZoB
zAfvXGnYjp5E0NJU6HLxevpGMdk7iBFfCeKcLAwsv37UNQaywOMQc7vv3WZQlHDykN1PatxQLn6ARD8GGEf79dE/9AlkhQCxlHIEcpNocnLKiCbRJr2HgYyrX3ljAm2I
N9vpW2hd7NSCbsU1vShy/eCZzQSwj1+dSEBwkQrRqb0qQdNgtnd4VWBHoVyrxvysR9rOMyldYtNAB7cWVzRcKN7YN+iWSI0zfA+1UPUf1bKq1ZzMI/Zob+dgiIqN8VcD
HmcEzAtP6wSVwuUCrOrzcCHFvNiqQi1T5MnwKL4z2nLDyVPFyT9mkESy/hN/zYLArZY+XdSkH4lY6omSSWNTV4GRuNuQw9mqEzrmAq2vIIrmjYZGTPpx5fHkDH12aeTG
onptsk/0Y/9ldbmfJSHFfWtiqFCy6uocqcJNEWo9YY01VhSrvClioX7Qj6NorwST+NzZYjl3+RZht0Pm6ZIdd1iiM/UPb8MeEeONk3N2ya+fomHeVEsb2MkpI9P0tcMH
rPfj45nsVrGnZjsRQVmdmNolzqmOu5tieMqUWjwcH8G6IK0TAA4T5TYQv0Y5GHGOXneGoQWAqZ2hEbcYCRGSEvUwqXBmY1DQcPWW+PIO/B/k6wUqAwgtuSBStD9GAe5/
s+rOB76DbYGn50lpAm8GwFSUyk5Y9QcJDUpAi+88uINfxD2QS7EmhakcnXZAOxCHYUYki6UZvXxxsNwbC1FTpI0+ysw/RPv5Xk8TRiyely020EBSHJHZ3yqXAuOamI0l
9kbNbbqj2du6gg2obdJ2eGxLbL2Q0ZFKW0FpFg7/1dSIYl/8pGFT4uC2KATOv0Re3ApB8BDdkUWfThOjI5LGG6ERmIwqKLYNHqdiR8HajS4Q8k9JinEAyQQWqr+Zjmt8
zds27SAkuyz6cmNxiEvCVx8qXYrWMJxivu9Lsthw7oJMHj0GSFokR6K0a1LIPHB0K/pH75N3B7NJmCypGGpRLcUoZmoW9PmpY6CoyEjD4zj9sAPGp/M4vLVk0ANIO+uP
mArLXJHXsI7Iwcf9ahqKFUNWpd2TShb7DPkitMjvdFCF+VUfJ58+FiJkLcaIEJPJiYwAh/bwVP5eS9N9xLfmDAS5qt6PiCgp4hsJjqU7f99reMrq4EsTKffdyBNRjHCd
GuhamFzN78+WfHL49mC6k7Khu5Fos/Svei9+Yt2ue0tSzUQfACadU4AiE9BR8llUnYX2AlynCo10Mt1AUBHwG3UTaGrmWxoH+fP/h/J4XxKFpTkeJHeyQGzsX4DaHyZ2
n0yu90p7+xGrM/MLzRymZViiM/UPb8MeEeONk3N2ya+fomHeVEsb2MkpI9P0tcMHRS9AICG48xoIeU1rHr11mNolzqmOu5tieMqUWjwcH8EEmAKBJ7Tzx4JqSEnRL875
XneGoQWAqZ2hEbcYCRGSEvUwqXBmY1DQcPWW+PIO/B98a5gOXOizz8CVLzw45O7Xs+rOB76DbYGn50lpAm8GwPDazMNb0znzVi5MyqK6dKBfxD2QS7EmhakcnXZAOxCH
YUYki6UZvXxxsNwbC1FTpFlYwCzuOQXLJx9B2jAEV3U20EBSHJHZ3yqXAuOamI0lCr60HrWqVthJD9K1t7euq2xLbL2Q0ZFKW0FpFg7/1dSjxtD53UgdWD9jCxxTRkkv
3ApB8BDdkUWfThOjI5LGG6ERmIwqKLYNHqdiR8HajS45G9829pAHRsAVT0ywk/rXzds27SAkuyz6cmNxiEvCV0GoAqpsHjC3YVMSJhlUtzpMHj0GSFokR6K0a1LIPHB0
K/pH75N3B7NJmCypGGpRLeZia5GeLJ+rXX5pCwuPaWT9sAPGp/M4vLVk0ANIO+uPdyyjfhGAlYErObiF2HVu9kNWpd2TShb7DPkitMjvdFC/D6wSZHzBU3jbhlbECgg6
iYwAh/bwVP5eS9N9xLfmDAS5qt6PiCgp4hsJjqU7f9+hBLwPSdMigsXIvHljeeJ6GuhamFzN78+WfHL49mC6kzBZRSUtUBUqspdfE/K8lxxSzUQfACadU4AiE9BR8llU
nYX2AlynCo10Mt1AUBHwG/gyAp7D8PKPNDT7WWVxdxeFpTkeJHeyQGzsX4DaHyZ2K5TivjNuJpbwi6O0qOC8fFiiM/UPb8MeEeONk3N2ya+fomHeVEsb2MkpI9P0tcMH
zn9Sb322k61bYwX5h/hMqtolzqmOu5tieMqUWjwcH8EGw3G/HBMe1YlvuHfEep44XneGoQWAqZ2hEbcYCRGSEvUwqXBmY1DQcPWW+PIO/B+YbjIGs+9XgyrZxvvF3ySi
s+rOB76DbYGn50lpAm8GwMtyXU/jXBpUdXtVehUNW4JfxD2QS7EmhakcnXZAOxCHYUYki6UZvXxxsNwbC1FTpA1w89ILoFWCRP9MQzQ+2f020EBSHJHZ3yqXAuOamI0l
AMPWcb3StwhbkSh9/AfTcmxLbL2Q0ZFKW0FpFg7/1dSmEMIFjkjWE2MhIcGr5Boz3ApB8BDdkUWfThOjI5LGG6ERmIwqKLYNHqdiR8HajS517j+Ai2qdujquViNqEcNw
zds27SAkuyz6cmNxiEvCV5TOlwYZ8EWQmRfcvXQq5LII5bMeKlQfdf9zZLUNMo/Rrk42U9mHCGJRqMPbIkkYB6e97lC9JyHQPiJa8L6IryXN2zbtICS7LPpyY3GIS8JX
U0gUP7XTUFAfcn5amVGbh5PMbmo30KKY7cjTYhfKXjUq1UpKHwPOYlYyPDYZ6Ib42mYL8x4PsvzEqDqGUPXUPK6XUDIMnJ36H9arRXPb8NzuAyLQfeXS761fW3yc9Wg4
TB49BkhaJEeitGtSyDxwdCv6R++TdwezSZgsqRhqUS3DWiPhdprXI899YYTDa9IChzJK+fRc8AUay6XSQfN19WTQyD6Q6aX0OqrRl7OdVqJwLvMRyoXMhTO9f3SLuPCR
bDnXjMPiOdR65htcTFryqPKdhQTe0sz1UxiGLzU/u2ZZX69N7nXKNEK5cxrpKBVqHT1OmfdOByz/DbI5/sfpia5RWRtLXpXkozZuEtV2KuEeHJwAezOKGDJrKAE0qNC7
/OEUtKYgPQdzI4gVajEb1/2wA8an8zi8tWTQA0g764+XrS1hOSrwtVxQPkcvI2ngFvISBihtfhwTEt+J4FJpqV+U1fs6V4PhGizug6soFAAWJwZ0Yt+2q5AcLEOK0cON
R9dAgAvBMrWvbBvhO3x839MPvf7u8TLeNqTuVwMZL+mIy8VcvpBTtqPuyToCvAqn5hLdV5VR/OWQ/obplGwvFAgTjI0okqjMNLyeO7Nc2eLGtNp9teJUOH9AqzyXTicd
hEKIFNbGkqH6Bv1RwghlyV784Jglm+S+QiMUHe51YdE7u9lNJoRX0KnYkwynTo1LaAMg4JXbEXHSTlqHPVHDWxwpACG5YtG38HqqHpXEnXmuh9YHHpDJGsM1cb5WM0In
BHs+ReqPckCgbOR3NQHRoA+0xpxRppEozxw/819/5mEH/ArauI/7JhlIcOQcaAsPc5cn9INVj8u29SDQMGLiii2Aipfj6kd4siAkaJNdYl0Ya4AFsiR42wl1/vo/t1kp
yVLDTH2mSf858HItLGLPExfg0VzntLa8CeT3kJ9sgsS10K50bkMhyjp2Benuc+Xw2Qy+LxrZxc4CyxDNOT7dim9WEWG9gV9Pzm550ouDOOofuqyez7d2uhs6v7M6pAhb
uOaeVhsxmWLryK4TpArsAXpZ0fXYYYRStOebRHoUJCt4CPW0l4tyy9p6yzBqgnjr6rc6Ji5BGTUXvf/h0ABIa4NCAjNU17Jiy9s0i2TUkHhnleZ44e5CJZiAmN3JkFRM
MNOOkhrq1r2yQEMLd1mxdO6u1BOQe0QORWI4AzKA27i/Wyba9sZ+x4wnpxI3EIYup15jCTU4MpepW/ksUw3rwlt6K7gBPJm99yV/QV2PBle1avMVhTtV/HcgkCZ6I/UQ
PpA5f78P5VnpcASrXxsBEzAoZ0QaXY6GzGqmJBL73Hx5w/uQMiCv42lZulpOOvcBC0Lc1hG7kZmVEIGpI2JPcJhaG+kpSAH+DPZDJwrX8PbdYfkNAyYqKkyNGSD1dTbY
yKPf7t4Tz4RqzMtLjVz97LQfdVXB1IPauf5SZKsWWgiTqK1r0PVuaNs56yGqb6VwCoY6G+aMcMTzd0Z2Is4/fa3iB18qAL+sPILzASEfU1YLQtzWEbuRmZUQgakjYk9w
bAXw2j3NH2z1FCTVsqueK9H2yl/8p0UkGbDWs6J5cbmTMsvt2CTMXHBSo1ak5+wlWVFSAhtzUlrSitIFqIXeXGldM3A8NENLO5iLQk3LAFWxfDfyoZuPQvJMtG5jQNxT
0w+9/u7xMt42pO5XAxkv6an2JmceLHenaqk2hD0+ZAbmEt1XlVH85ZD+humUbC8UCBOMjSiSqMw0vJ47s1zZ4ut5A3JUcnEMaVuDl7fLAJSEQogU1saSofoG/VHCCGXJ
wUPqD2dolVh8R9w9pcbfrQsH6EC0YTBY4Y7QKFjezw9oAyDgldsRcdJOWoc9UcNbOGTs+WjqtSL9+6h9YSWg4q6H1gcekMkawzVxvlYzQicEez5F6o9yQKBs5Hc1AdGg
LxZ1G+tWnuEWh9SoDzkX3Qf8Ctq4j/smGUhw5BxoCw+6L2SRvbVtAV/tUMqkMZCnLYCKl+PqR3iyICRok11iXRhrgAWyJHjbCXX++j+3WSndN6ZiymzIWp7eWteE6SKy
F+DRXOe0trwJ5PeQn2yCxFcfsrQtsp8FZ33chkiGiqN3N8cusuNUsYNKmUBpywgmb1YRYb2BX0/ObnnSi4M46h+6rJ7Pt3a6Gzq/szqkCFvN2FzQhG4LtmWyZosAd28x
elnR9dhhhFK055tEehQkK9DiMuF1xp0ZaXqOt3vzzanqtzomLkEZNRe9/+HQAEhrg0ICM1TXsmLL2zSLZNSQeCVM9LiXydU9zbK9+d4eclkw046SGurWvbJAQwt3WbF0
RSttSCqZzDqpfyee1VOS8b9bJtr2xn7HjCenEjcQhi51+YWr2kPkI5j7Zaiity+guHgZFS4QulVBPqMufyEbK7Vq8xWFO1X8dyCQJnoj9RA+kDl/vw/lWelwBKtfGwET
2W3knJB5OR+PgL+aNaYZjHnD+5AyIK/jaVm6Wk469wFns6vWvlHyc6/YPo9HfGS+mFob6SlIAf4M9kMnCtfw9t1h+Q0DJioqTI0ZIPV1NthOGIrQ8VZ/PjxHpONjsV2i
tB91VcHUg9q5/lJkqxZaCJOorWvQ9W5o2znrIapvpXAGKV4R/aSNu0XWFzEsBVzg7XGZ85IUQmW562sZyLhBEmezq9a+UfJzr9g+j0d8ZL5sBfDaPc0fbPUUJNWyq54r
0fbKX/ynRSQZsNazonlxuTu5q4QHK7UsKOrQaLck1TpZUVICG3NSWtKK0gWohd5caV0zcDw0Q0s7mItCTcsAVc0SIWBPmg501lkQfcEocvzTD73+7vEy3jak7lcDGS/p
HCx8WGS3/JYLKC9Xdcrj3uYS3VeVUfzlkP6G6ZRsLxQIE4yNKJKozDS8njuzXNni2mHYjZj+dWwT9jxNKMzLfYRCiBTWxpKh+gb9UcIIZcnGN8EW6KXHE+6tt/7XYvlS
jMlCGIACqJAu9ao2fjaZU2gDIOCV2xFx0k5ahz1Rw1vlfzop0d8ZBq5vi91Kg9fcrofWBx6QyRrDNXG+VjNCJwR7PkXqj3JAoGzkdzUB0aBH1yOn48e3WamOZpSRkl7q
B/wK2riP+yYZSHDkHGgLD8dgGGICar/mlgS2EKZqgnwtgIqX4+pHeLIgJGiTXWJdGGuABbIkeNsJdf76P7dZKbpfmFVnagUa977M2ieacZoX4NFc57S2vAnk95CfbILE
uooWJwln06p12vIduiPyAHMq/D6dwQE3PcVY2UD48rlvVhFhvYFfT85uedKLgzjqH7qsns+3drobOr+zOqQIW2wfcYQ2LBMqi7aJ/SsYLO16WdH12GGEUrTnm0R6FCQr
4bM6r8O4fsR2A12IpDiD56Nc7lQfOr8UC67djcGj/1exLJToS4d3h5hJ/sWUhKhTHHLlZ1BhwQpPSmMPn8YykAFgV5qwBQBy8ENOub5gORwfuqyez7d2uhs6v7M6pAhb
k1hqb2TtXqhtuN85dPF15FYtBOGCz2zg05dbO4rRtPVzlyf0g1WPy7b1INAwYuKK4onBMNfnj2OSdWPIOZzKWludtk+PC+zxOsaSkSrCRV0U5OQK2mrVyCJgjwA6gd2n
k204EKx0tCOl3v6ZmxOxiMKj8OQiS2FFlkSpJs14bu8TVbYrQfC1M2qYLojD7B7f1pYzMtsKf+k3TtHXiFO5eFLsGTS4q/MxNXv3ibenpNotgIqX4+pHeLIgJGiTXWJd
GGuABbIkeNsJdf76P7dZKeZ6RKGaE3ofNlEzPQbTmqEV3Ck/hipa9CMZRTN5BsJ7/Jkb4QHkR2iQ6hX0/polyO2+qdlYEE61541/ZIzh9MEmJxHUH62HdYaYRttFVx3s
tTVcIrU/r3vvRt/AWM+B7ClgA3fnaMeY311QRMvWBSJ5w/uQMiCv42lZulpOOvcBc5cn9INVj8u29SDQMGLiiveWXmtVqBOshG2tfzPLyXQYSbjrJSWBvl0YVCndIMpa
POk+4k3gLH8UFE/IzG2FY5hHvulE7ei5xUHtUepR0jg2hfbdEQjGXg8MLLAyfRsPiYu8xX3qSyoCp7gTHIYz6P8jNqhSaTlVFp5SNs8CWWIWZXlyLa64DUSH7bWvFcvv
NbrcaOgcHGrQwaPOtTYJK8+xRhjpnGbNY+ZkusHUtuSv9UWhXRxL9r9N2y9eEF1nQZ1LKj8lLRALMGvwgkmcesbVSmGiLzig9VyU8IbhHd2t7vyqk5BM6riMnHax74HI
ob9JBPK7iGGksr+a77v3RjFwnm49aGXc5rxcjLmBS2zuKCL9Lp4g7UMjGHUs+wFxa61JvRVhBE9bmdSU3zVH5I5yhuQdhu+zAi6TOkOi9In74H2WsNpUNWxKT9/nwKFa
+iwjS5jbQFDWrXzj1HfGWT4jfJhENGsE243u+iag7hVh7gw/+V/xENi7o9EIviJYZx0zmJETrVPJe5rPUD6Amek6ixtg+ulYgU71fXImZD2seCbIBdkuIoLdYGxBqhda
6VHtcH7Qh55fItyo2eyYsps4nP9JEH1oIaDJJ3KwJqWS8h+VhbfFlExiul1Jzs9Joe9hNfqRSVhGx/RpsFYJlHbYaUg9+J4fxNek+YBxVyu5E5e8tJwuUeA2bIpqYFIb
wbyUxsmQPkSW+sZhnDZ+KrTWEowasSMj3VOsd+ofNUCAWnW6xewiSSozewz7NlDmE+z0IFUBtcZE4frt0KRxB3CnRlQDUok9JoHV2LZCyxfo9BjT7V6Jrt0AllVzRTiz
IRMkBLNBT8E7VfcDsUf24v/W5TQsGpAamw60G6jUis7Sk7/3RFROdUlXuuimyJFgWs35EbY7/qTBB4LDozjncDthk+t3SyQjLMHjntBU8AuqwxqdP2es+1NAVM7eEVOH
TyGVGl54tAj9tpHT573OO3Elo5sZt5bFFTs8gX4Y1rpoXFJMT7YwKAx+S4D3XUNbhDF7vI1gWAb3+zvUrmXXCN+v65sPTOXmj670Iu5j/j4X2z+7RpLg0q3aMMHrLnTC
Uginsy3TpVneOxg9th1Tec9NGq5Qi7I9P9RnALQ5CsMmVDiUfzVOeLTcKB3RTHpJuoaCvUBpl0LOZAYd738IJHN6MIBX1pV9+a1Gv3V4fkZ8+ngNTyzkkvV9fTjm9X3M
jXME+RMUZidKNgjPXTJrUMvsCSqtDb6KNdIYFmrgDXbgtmfxn8ZAK8cmNUY9Arc7ap9z3zMw1QKVUntlZ8KBHLXdMCuP/Kow53tSE02Ypo7pZ1xgPSj5z0NsMgV5RCwb
lYou3u54ygT9s+OZQ8fuN7BJJXjXuVABDQE08X9ysuNrjkBAT4K9Fu0Qt/XM+emiBOy/vYkUsiMLeh+ilqKeLRrgYDkJAgXt4cQlk1/alW3NuP0z48ciqlON4BmWHtEn
DvgCtnewHaBZT2SdVjP3zQ2gsUZ+ctqxBxL/aTMmaotTz0sQXH3MVbtV3cZz0HlKbNjDRcvwE1BoGvPnyFRj2PmJBPFab9sxTnVJR1xte+u5YoYDbU2l2IIyNSpVPuiy
Mm2g0d/DuowWzXfdC2XW89sQws340GaeJMAHLzfWw/Vh1PpizIHCvbB3w691ahiP/ljQisGm20MyY8foiR8+aFEARl0IGTqTiVRPWzBqmztaOWrVapR9/Ig2WshrWNNK
99ZU9Id4KkYj+jnRS1WcqQbyXVq0sQ0Ufplt8vwtf3O/53cCmI5xcjK3kYi2LJwVuWKGA21NpdiCMjUqVT7osoxVGCG067by/Yfh00HBxYQAPM4tEjK7iYsN5uMLgI38
sUxehEhMS/LGLCtCN/KV7ZcYQURHT00uizYO1XhCtaRYBfRpKryN0+d9ih+Ddagdr0QmjCn2/KtuskejV8wFH3PVDwTXVZ2WxfAT5ReXKFRdKOwO7G+90uDK6byk11xP
0gu+0siZgpup1A2MoJfBZcu6bpf0koypEhaaTKQKyZxRxzcR2Yl7vEleYWs/4cBS9T5CMBCjEFDbLp5ze6ESBeUeOF8/q08ndL8bakTwWZGTTd9zo9gXac2imlfVhkL9
fIc+LFYiABY4ZQF5z855mAXisuskWIqjlpGSn6bYTY24BJXQ70QUa0+puF/S4lgleednrdt/LyamiZGxjLCYBQMP4l+DqRuJJ+dDXroTx2dzdSSz5S/kKQmD65Oint//
+y7PldAGP9Um7NPE5IiWFk8iUDKGm8k2hmfx3N+Mve81YRfqmbbOx2Y0ynYgGFeU2OQFJmi+WpHEvJJYCXSZC5CJ5JE+YPF02xH1LbNuUCqVuEKZGYuAR2xEG73At4Tf
3Z+tShOpUa4tEKmlevx/vNbT8G4dKx7Kl9vKy0/jrSc92l+uIF6cxJYrV8aFhivMt9HwYtgZp4jdJWgOmT6r8UcuQWL8VUWKOqV9t0cIJdfuWMg+pnd4mpXUPbDf5Wbi
IdzUELr6OGN8CA5vDjFYUYIn1rVNId4cRcwiJViwTj2dzGHJsZubjUhcLL+3a5PDOz4VyjAcg9Zlj+cwFwFDXkw6J01tlUWWFY0eaAd+0SV4FUbdERsxVUBipngBOGqC
HQ87wozU++4tjaY5ADzpvPRUN0EwXRZZn7SuhCUQi9ok8Ks9+UX76NA03Bw7NDhCIjE1GaB+QnvN5t/w7sK8ymTJpIwpxkycGRJsy7JdEubDwhaZLSo9wlHlDop3iHwv
gFKh0E2u4dtRh+pZ+S3e3kw6J01tlUWWFY0eaAd+0SWApjcc4q02He313LOLF1SEEIks5L4eRsP696OBQBRhwQx2kKBOqdgyqGKhGKOdf055OlaeQz172pFL5baV0Fpt
E9o/JX5YGXcfm8vew3oPnyLlg5xiMS3smrZHHY545/VMjBb9uMviGDlQiMLaZjgq6OTVdnE2FyDiiztZEhE9ulDhScGQMisBMGbux7SOpXz5PbD0RDaxZu7+XkzhLnoE
mA/1nVNH0BKbY/LPFewctGzU8kIXWdoVqTtHfm13mA8cWdHPYxB18uMkj1Emgh2F1egA9uW1ApoQehKqnVM2LeZHedJVs5+VmpVNLPesu4OAUqHQTa7h21GH6ln5Ld7e
TDonTW2VRZYVjR5oB37RJQ7f6diZ6LcPrbzrI1dj4T1fiM8bAmEjRVbNz06Josu1kJe0dRu9ydSsdAOeehmyjhy44BanweVwzVmIOYH3oa1Ppn9l5Aw4aC52FIsRpNYK
GAAhuM2Ni9ofyDfTayGPLogWwAkK+/H9qs1RP6cAm0Nkjb7owkbC60XvVJHOWzyUDnEB/4fVwQVRUgJEow3qsjFsUnBTzIxtGAgPeKk80tHB51hOD63lnzcz5x7X2MCu
yM98aw7QKE72KX8jppWsBU8iUDKGm8k2hmfx3N+Mve/K77RB6IEtqVOQ2ENBHstxeOrlEqKdGKAqDcSRP2GkN8c40kxf+lZn34bO1gpWUTtjRiGeRZMxqBXBd/ooD2Ty
wBzToZTWGP1y/HEvRxdUiv51hvbsmYwWIcJyUB1xMhYj+Oiii3Ru+r5VVAzj0K4g0t/cDwMUwJChx+VfwTfoH3hQyz6U4cnsp146chnJPwipke42a8avDa8r8kKYOYu9
KfM5aJKCnAkf+YQGKz1q3G5ptiiUWrTIqDlYvrrlvczv4iUpwckK32ZLz75pBe5wm9gTYeeU0JPm/IMCBezRaRxOrdXUxq0mJ4K+s7B72YvEa3Q+d9dwWEhkY/ej/6jQ
ZOfDb0YOZlyjO4u7mVZnNgFPEUlqloXxqUFwoeqdSThoJ7QVKM84VlYWIwJEpo2eG2Zetz7EzdnQ+XE5H3mDN/lPUeZMNeSiOMuTPb39mhIwNIPSfpGUy1T1JaUzhob6
UOFJwZAyKwEwZu7HtI6lfBiQioVVj6lgLGOCqVcFvaiDn104E3+5tRITT8ciLMuuXxL3j1TkyvfddkNO7uD1nTDvFbO3+L6gpZDZ5IjvnS/EYjvMZFCsfeIQrq0rbG6j
tWtHCQAgMoQr42sPKIcpFsSYE9KTQoJnkpNUEuMBl4G0txuXfEcFVfKM1t8zie/TWSqk9BNcixaZ3y6e7wbjqx6YK7ZBGPRyMzt2FhZ4swsGHU8gh+Jkdb78oFLSoqWZ
d4ocn89J25H9Hepme55/xSP46KKLdG76vlVUDOPQriBwqVrkfXbwJ52w+OLaRpnXW6Z02B7BRwwANoZYiOj2dCIR3P5p4AEH6GIH2mcqsM1Q4UnBkDIrATBm7se0jqV8
GJCKhVWPqWAsY4KpVwW9qIOfXTgTf7m1EhNPxyIsy67uSMc9kGMS6EzcRvGvYkCQHQ87wozU++4tjaY5ADzpvNHsB8rczOQMzu1Q5+kHNDEMyDtUDOhZkWlzK1RD8z8Q
fIc+LFYiABY4ZQF5z855mBUEzBliB6w6ekqAAXH+OzTrvYkqeoX0rTLCcYR8ld7VkJe0dRu9ydSsdAOeehmyjhq48TVXgUi1cnsNxpQayY3bEMLN+NBmniTABy831sP1
xD4dj6qtCVf/oHiMMOjruCbjIKhhvpMgVz1f1e+NNnIv6KlKHFxHvDex2lVkN3K80d+6ncxwP2/SN8en/135vi/r/Vx2xS7f8cXo2mKf6rl9/olsnwicC9qc5eyKNIHr
pXKHsJV0YqrkbXM/od8iOgwj2EnwkTs0LkvKPNNFHozI5lam4UvfsoAoOMUpGUiUWAX0aSq8jdPnfYofg3WoHRIkdoA29Hf8uAo0+z04f4pR2c0+AkWAxu4CN+/n6D87
t50h3YbP+u9syWuxY4+VmgosB4ctwpUJhSA5jW7vtJL5A5olJ/s9qkjzNcl90mLA6t9Kl6lhXumSIyrGIibuBZ5haPN3PCGs0MVjW3HenbxJuxLwylvCxGynszkPlAjs
kFTXiwrzVXLPni0aEIC4PM3OqvbosFkAM/spQ1QrRbJUAT75dMSsuhE1zCmTvZgRxJgT0pNCgmeSk1QS4wGXgXjq5RKinRigKg3EkT9hpDeK4d0aMTe3cwGq7q5Z7M6C
NTpfnag3BoKoe8AusaIomznupGqaHE11+ctL5I17EHL4QYBSObw1rGd3sXA29GJVW2ufW/6Fc7g1WJ1W2zvjWqL+8sBAYnDeYAF5dFVjshIVrm6DuZgUttkjwiXLZ41P
iqufVS6TOUhCNpjOJbgnTm6KrJlHhzbSxI+D1/Q2fd7Fdlo+lvK7RA19E/e2RvEU5eF9b1yPGe80Gr3rtI1eEOKvwfDvNMfswJomrSPIH4Y4XaLbxzNx5fD3BpaHiHO1
FNsNKqLTvOhKVi2GlT8QHZcYQURHT00uizYO1XhCtaQQiSzkvh5Gw/r3o4FAFGHBr0QmjCn2/KtuskejV8wFH0L0gP8gcvMpiCB+jNz/IZuBs/aMd8/B1/6N15driCId
Oe6kapocTXX5y0vkjXsQcvhBgFI5vDWsZ3excDb0YlVXE3UUzBFTw/0Ehr9cC55ddJuBBBvZlSde3VhOTgDmf+9KNMsRDRUdiCGeqArnASSYdz/ucvywc2SsG9P7kIZM
fphmSvaqgov8aJB+sQ3X/bLnWBU5V6OXD0OPG5TfD63IpZLopKlgAOuv1gikzXeuHQ87wozU++4tjaY5ADzpvLVhWHDNbYLLZP7+SRM4eRKmp9epKmGNBRmlJmMfjKB9
0gu+0siZgpup1A2MoJfBZTmM8Cfr6oT+3K8zVcs/EnZGE8nML2v6dHlcvAYEcAxs0t/cDwMUwJChx+VfwTfoH7LnWBU5V6OXD0OPG5TfD61qBR17tWQpht24Vd8GxHAh
36pfX4Ld3/KDRRr+7E78ueEn8a2nOmEQQUvLv/ScFn0oGmIwTJAunkLIdFY6HGeNm5h6mxfQ+nbo6TJvjOC23aIH56/mN+Of/D2XL9C2XPRL0qPfvLuLpw3E7fNczYFl
XZywK2QXd/U/gcZGStaVbGWMr17BpgTVgEh6ikJyP84YACG4zY2L2h/IN9NrIY8uEzMNm7fCBdYuIMlQTJtn02SNvujCRsLrRe9Ukc5bPJQuhyOrGQtPuxiqUHn9x7Zd
CwHGsRWqqSXEBapUE4SMi5Ul2fJT8Ot7wRMN2b+G/5vj1keccCv5qbp+KlMxu307D5H2JYICjyhMaLWvx4yHM9Hfup3McD9v0jfHp/9d+b7/1DTjvJEeaRwtrHvx8Hno
g58RaUrKPR787K+Qk/hj66iUZUq0r/px5W+qQYIyYFWpuNzDqhLsWuUV4zGQ7UE7/ljQisGm20MyY8foiR8+aL4GgqxyOJLuudVrtfg9gipaOWrVapR9/Ig2WshrWNNK
erwG2QImcCjKNPXZzev1y0CcsebCkn5jiSiOG0cvcZWdY3Xu3NZ9T9TYAh7WyFhR4+XQbul+MF2+3rH/WPkKAeKMmvcPbVr1uChz/GSj7/Lww/YE/oTw+Jc3rIDXU262
4Sfxrac6YRBBS8u/9JwWfacFH16P5Y5mFCCMf0KJGxA92l+uIF6cxJYrV8aFhivMUseiV5sNdsiV3Gc/myEE1Q24jrIlES4j0PSMaJufZ5pS91hQKYMUxip5sO+MhK18
qJRlSrSv+nHlb6pBgjJgVam43MOqEuxa5RXjMZDtQTvxq554Ombp9EdvWafZiti/hk6MOHFi3sMVWRQgKURHFYsnZXY+8KIQYQ74qqtSm1DngcF31XJvkjW/Kwo5s4Xg
EIks5L4eRsP696OBQBRhwSOoV01L7+igawnbk4+zTYaVolUHfLkCdd8RL4ADgSEKdJuBBBvZlSde3VhOTgDmfzJkU0HPt2s4PMAVb6E8wEZ994YFWdQQaC6qVtmWPcwX
F3N2vIhQOOY+cHZuVJ7r9UtXviK4g+hgI5STUOwE1Y1kSSWOK5OyJ0f3cKOFeykQWAX0aSq8jdPnfYofg3WoHRIkdoA29Hf8uAo0+z04f4rcvROUB8KxZE5pDSMrcup4
RsOzWglWcbmpGWCgnZtvVrRqHduNBYNLr/jm3OV6nsOSMVmXvUU81b5kO8UbLu2XokttMty9uDO4VHZ9Zl1m33uTbH+Vl+axKU5pa0FoxfmUNa0ehO5G+f/K/Jt/nsXM
qpmqWKdJ9xKIn4qYuvwJbCjIpquihNjFUL3UXN6ORG/J2yL9tPwxHYQdi0jpq3Z01iRbfwI+9T1KqWhuV2gQ9C5ikYiNpSLu1/ezzjFq4+t4MoPh6dm90XZX1jegsSbJ
NtXnXeVzf94QRinks/40EZkjywgsMW+sqR1fT6+IfxuLkil0UJwP4VVNvOw1v37ZMP+6O3G2HLKuETV3FrUD3oGBLFyt5+O3xxf8V6ZgzrMdsngB4V2+oYR7XaXeD8Uc
wcBPkziYxASvode8/amCWH/et7dxOR+Cnjr9Unfo7PLVYSZ4BRdgtDOinXALiMASCkDWMJYo66cNRFZO7Ne9GLZv2c35Zaz8vKDhVR1NwbGBgSxcrefjt8cX/FemYM6z
23wJ2jDRjEXxrTJWMzuOOyt/Ey20GxC/mihrIsICNcoNPYo6uxP2CPH3Cj26adE/+omNJdwT0mz7NiIpTqfDfQpA1jCWKOunDURWTuzXvRhLwVd7b6HTQSA5hwOxJqyM
W+lrGvIKcN0xnddeMOy+6mdrC939cxRK7NSZzBYjBjJIRW47wBeiq//2+FWo2DSjrOfNHGHYnsD6y55PZYYTdT2u5hk0Qpg12dl3+TlBb3UsZPf+XUbDRE87OkAkC999
3tg36JZIjTN8D7VQ9R/VsgXvM14FwxFYb1YqzjzEJ9RHbE8R0jHvFGkRAPbPyPGB30xkJlUwHNVlgYCWv0vgYePYpK9igx5sBhjqKI3uvc85Qn/kikJsIju93FX3s+qS
bJHjTpMSi9vK8j5WEMQwx62WPl3UpB+JWOqJkkljU1dnVoxou/InaFvbl4W1S40/Pa7mGTRCmDXZ2Xf5OUFvda6fKHU/nVM7jvaXG1y1K6HmjYZGTPpx5fHkDH12aeTG
geUE7x5eBm0ilUw0a1vG2aLlc3AAD/JPSPlSGakhd0dIRW47wBeiq//2+FWo2DSjJCf47/tWUtIZk8B+Fqpr58qIJtEmvYeBjKtfeWMCbYiIHtA50WlszBhM4/y7s97N
NtXnXeVzf94QRinks/40Ede96NSCkQoVyOyz/7cf1t3nA6fPaUxFqBAd4MoExW1NY3pLPGnMEHj8qazZADYd8obk6UyHe7aiBUOb5S6hWPk9ruYZNEKYNdnZd/k5QW91
hnyxrYgYrwzJp7U0Vtw38K2WPl3UpB+JWOqJkkljU1cQsVbfk8+7MQ+REEGyIII6pxk+/GuInDR1zAlboPqOnmN6SzxpzBB4/Kms2QA2HfKc1qtaXyuYDdjLzQTYxHgu
4h49K08aGem0bm/AE6/r5sVm0pbXmQjWooa5jiuDxD+6ASOCW/GjBkbjl+btxHNq1OZJ0M8rBGRm3cio3yfcii5zNzklqzTDF2OUaKTP4gjB8NsHEAay1aSm0UtDBQUh
qjLUzPoJ3UFIUE4aFqAvrwHiDdnMU4+TqlYmhDiSciQnIvsyOcqpLLK4U2cDdSEgz4luRg03VQnxFTCF9XkLDfKKhBsoiKz5v2LfJG3/NHBM4x1hVrUC73d5DN/0niLC
DuZST9OIBBbN7BdsMC0NXyCaOm17/GtoJRxqT7+J7Z/e2DfolkiNM3wPtVD1H9Wyi/OxW6RoZro3XIf5QSmptR5nBMwLT+sElcLlAqzq83DLtxKF8BX8MTWfIP/0yon3
2LnLEJ2BbTShGAJXavcWUvU9TpKRqZDWXuxY4ZfCwnp2PcIE0bAIKuIWvN0AnLVpoWWJOiwPCsTVlp8tcMkZWft5gkSMMrQVtv5RLHuP67kgvXseuPgL5fysh2hy81Qi
Vjw4aXuCnsavEJ8bfn0aY+v8dCuUio3DyNTRRCnDyRkiacOQPNtNa20y9f0ZdYpHWaFzyF99kpePBbWVPNrbEqzZ7sY66qLFgF6/MgCMyfI7d6j50fh5BIAAC6E5x73D
jDeRlaIBVXZH/++wOpd/vVY8OGl7gp7GrxCfG359GmNhYRjXEmSvqAKVR4PmkrrWnVghlUeBzK7WTo2AcEi8szO0tTYtrCrLBGjQSAgZvOP1C2LpANfl7PGh5Cto2yEv
T4BBo+2L/jNzjFsVHIKffsXTavLQIltphKVE6GDEgFyzISEHY+kgJNRUkJcfcWjvbEpWVUfh4NbUCHVH+8Jg7gxaF0j2FyE4wRcHqOkV6ni1X4HgfkvE/AK9GJUblTb9
GuhamFzN78+WfHL49mC6k1pXaqwjTWmu+dqwWtwYflFIQT9EhQ8z+4rL4XsDkE0hN8RlU4qQCxVAnzTtmSZc2WNugVt2dbz+I0O0NVi7ZujC3/00FfeX3JnhsDCNOBnj
q+GlZ2A93HBvhFgkDA7XU4uObAltXSZVBbfUzGUweX0x21lGxClIQPtPprYALnYxCmWl0y7TySDsue0Kn8wCIJJ55xpYezQTAgl4bs+CYN6N6Bl9lqCHJdyAss5qoda+
qXghEQ7eaItwNKIaFBqiwJ0bvupPSkv/bkE9dD0OoHJ+AwS1qfRXP18pgMdfiQWFIBt6IBH7qcXdWaCiQbbWZEFbh2nsIeENS5+vei/Hqo55lRZlrYe60rLWzYWMKxV6
BK9hANO2+eDDVECkBPZwWi/r/Vx2xS7f8cXo2mKf6rmXbN/It7wAITwXoyEL/vJJErXOmxfdForEPQLIfFSOfZvGSSV0HGuNfqRWiVfsjGfDAVEi4t0nOrEe04ujexFn
bEtsvZDRkUpbQWkWDv/V1EtE8MzCYRDLOfRT7cHQjDYD/WxJpu6bRrn4hDsIxZNK5zbe2d1YIJhmBuZnAg6erGCYhPLpcqKju0MMDRKgZXusocuO010WhyqyL5G2n15O
O0BUPmRGPkRlEkutajL5UUYFzFeWPAkCePtf9EFFkdNsSlZVR+Hg1tQIdUf7wmDuDFoXSPYXITjBFweo6RXqeBl3yYh2FfpW88HKe4V+Yf8a6FqYXM3vz5Z8cvj2YLqT
4g2+fmVs2UZqqhCH2jtWBkhBP0SFDzP7isvhewOQTSE3xGVTipALFUCfNO2ZJlzZY26BW3Z1vP4jQ7Q1WLtm6IivFo3sxJK5y+E6lsKqsY+r4aVnYD3ccG+EWCQMDtdT
i45sCW1dJlUFt9TMZTB5fcOhFeOnkHPV1T/h8BUmHBUKZaXTLtPJIOy57QqfzAIgknnnGlh7NBMCCXhuz4Jg3kvSo9+8u4unDcTt81zNgWWpeCERDt5oi3A0ohoUGqLA
nRu+6k9KS/9uQT10PQ6gcsdMQvWKoXhU+7ag+4xvXg/8CvFL9nXrqXZvAioIb0/7AuV6qTJABMBBI/DZo/tVtPl3iKxxdvScCXKXzRxAdh3+y8NtM8KqvO1qX5gRUhYZ
/rfzN8nxcfJxYGr+BiSwLwYrBWcuJ8sazxAZfhUyIr/N2zbtICS7LPpyY3GIS8JXul0g+F2dtIFI3SE2tDsgvmoFHXu1ZCmG3bhV3wbEcCF5EUO3T6jLTbRha4/ORNC1
+mwq6GUFZ1E2i+vK+NiyJeO9q3mE0lrtIWzcUJCE6tBed4ahBYCpnaERtxgJEZISPv7KKydOb5DumOIYJ0rnmty9E5QHwrFkTmkNIyty6nhr65HkpVnEXVXyTEHELp8i
YgSKxTItS3FnWW19ZJdu3CWILXy6pwurX2swL9A2HdFe6h/XczmMHOQv/fCjUDooDGGjYSX/mJhUZdMFPwZj1uD0WiELlmxbonBLzT+bSKUjjIGU8fPjpTG7l+GfYOCB
r2piFXVQkpq3Ns49t5xos44LzwAFl/1TNGWdpRt0dRdEwmKjJmxNSGuZCY4zmuenNw58zosXOvPD95MdEF7hW+1kZn8UwSFaPkMSTtF3IQSA25uI/3gl4cSEoQKykgVG
s2KrrT5cUppAsc2lxf37ltxqvflzjvx93bNY/C+gxnCCJ9a1TSHeHEXMIiVYsE49ozhWY5wxSULmrmqS3G89vxpFyYDcBRXZ29WxDYkdoig8QDsuszWDXbr8+bC2UdGm
uUz8fWh3LZfRF8UJ+BepqO6u1BOQe0QORWI4AzKA27g/7DVBacZWp88Hr/bRDFRJOVx++kRPkQbMJK9Dx5Khe0L0gP8gcvMpiCB+jNz/IZuUBlFUdZ+OUvhHJ8nKwB6v
MoA6GBaA9uQBG/ZusBM7iuemef9cHGL3a+ZQlj21HV/l4X1vXI8Z7zQaveu0jV4QfgINDVETYvHoVQPtC3j14Qxho2El/5iYVGXTBT8GY9bv5rvXd5d+NFLqme8dJbGR
qXJ6eSD6pj2VLdWh3mrFXwrwCIojb2bMKlbuMAO6+LDoirqX1swMjGDL7dvFTAXbr2Oja9OH5WteH1G+nrZlqSM+VMlz5oTs9LOu6rO0XGbDP85JnttkNzt/lR6616CA
ZpVM+5OsccqDcGsxoFDShP3vaj7+R2ADfpxibI7Ia7XbJWwG38hkfHu6ChLNQa9ckEhE+JscsAzzIEdqIdzL7qNPaccxuN6y7QB6S5HFrFCKMqKODz171NHa8A9xg8iq
uw5iZ7eHFRxHYhSOqwj/8JBIRPibHLAM8yBHaiHcy+4jjBO+2FUX4BOvmr+ko2jmc9UPBNdVnZbF8BPlF5coVGOVjPNvuYMnO2hb7JwUKzaQSET4mxywDPMgR2oh3Mvu
fh/nGdLDRp7Bq4foHVSE9Mu6bpf0koypEhaaTKQKyZy3wW74rcm58uRZVRmNgKYKCG259C+NnaYyMaaa45ZUqm1pQje7mP7fRMkctRTcXCjcFgADc27QExe1nrTbzq4a
G5cCALOMDQ+cisT/xqxXjWqQvNHZBmeprRVFoOZcmMmbCCQDVrZwvpG0Wo4vWEe39gVqZU5+4yFzrjkX5I3mZ3BDoAs4+aT2bJkmAo8F0rWmTlfgDYiUHNOrqecYUih1
jFOM9WnaoHUzZQ9pHilGHtR/34D9WpARq3YX0WYzbe+4v8R4QN6Yc43syrWYdujgWoEgjlNIHcqeS5V1wqTOB+mgV4EUQRg+3ragSpCGf4Ww27DseU4sD37CTI6D63v5
CGBKdpFgtb7tT6EtoxjsHqnyR404XA2CpuZcm0zWBISXAySGzG9ewOhmMx6IK0K8gisfbmhDGQYqJf6jwlMGjhds7iCdd+imO2cPgXFQKSh3ihyfz0nbkf0d6mZ7nn/F
x0EajygqHKu1LNxnvdFb5jOUK96rS8xB48ZjyRZy2f+4/1n6FKlRVfdI000DfmeIB798itdKziy5/HWA0xqBYICmNxzirTYd7fXcs4sXVIToirqX1swMjGDL7dvFTAXb
Gr4R8BntroPbk7kiqCzsNnOXJ/SDVY/LtvUg0DBi4opLbYTiCDt8iUfqA2gWgnQya/58hQYl3ACOQcN6kTFx/oqrn1UukzlIQjaYziW4J04Q8t9DjQKIez/y6TbJza2s
huoFl7/sPZmT//qF+/ugAjrVzWI1oz0pt9FVebxAzPXLum6X9JKMqRIWmkykCsmckVDbADVAlhKdnJt85pdMBNsy7DskuCsd5dCC3QqRWLaXtneJiDh3sQPuF0HFHLP3
M5Qr3qtLzEHjxmPJFnLZ//503FIPftV/+iFcCbjubPPbMuw7JLgrHeXQgt0KkVi2Ndg7Sl9U+HdABcSeZvHBxTOUK96rS8xB48ZjyRZy2f8U0tFJPseXygklEunBjD11
2zLsOyS4Kx3l0ILdCpFYtgaMrZyQJZIQFGiR71ov40a0U5GbQuPLHE98uUjgU8otqXghEQ7eaItwNKIaFBqiwC0Uay10xBoFf0RJHcBpcaH9f2Qj3eYgdL/v3efXdFJS
UdopMJfETwJ6MKgXpP2UwIqrn1UukzlIQjaYziW4J060jQYu/kAO7xV8qO4Dv8pTWTA8N86wIl2HZajD3Qahb/ray+v+YroLAZagdzQ1dk7Q6V7BZXW7Z1BN6NEZirI7
MM06zAsD2tJ1Gn4dkASwNmDs1MJPZSJwLaqcbNbboj7NBUbW/JDe38nBUvFZuxts0wI4OQtVmUKfZC3sXS7t3QpmwEWQNASjWfFvDUORhAt+Cb5leuXTv2ahyIvuR3on
0kPJTQbGwWLbIFRQ6WbC4EG2eeINdbzW+yKWkPnh+6yLGtlDeTcyavaXa4wXxMZ57ZQrWY56AXQEAZqDhRp9glGd4g3eQQAh3ESq9YMdaza4N3qiJhdBNSJVksonmQsr
9FQ3QTBdFlmftK6EJRCL2pgz1S7+DXUK9QVv3ED+yHxJEwPqAxo7A2yl4zTg1I/zZEkljiuTsidH93CjhXspEOiKupfWzAyMYMvt28VMBdtL4L2PBHfUHgQXHFerQY2M
KlbvoBPNRUZX4FcODJke8EINjqSk8+jzkcHX3yn5PVW/liGvHepGd27YLJf10F8N/ljQisGm20MyY8foiR8+aMBO3K8sG9l7IOZZRpKQM7hKITSbTYJw1RHvwvS2sFVE
eANR1aLCvnJ7lVF+nC+Yz/fWVPSHeCpGI/o50UtVnKlvaiGtT0xI1Dh90dbsBlyXTkYHIcy3TC8KVrTsEavUFVrUQJzqEdfc8juTcDcewh1AEOY24sIkYsZTL8wivJJE
1TgnJKlSGCm7gW7awPYhmzMibtB2pQzFN3wighXVA06XGEFER09NLos2DtV4QrWk6Iq6l9bMDIxgy+3bxUwF24Q+ac2JI1VCjd/9nEcZJgQzIm7QdqUMxTd8IoIV1QNO
tNkE1Xbxwdl6RBye7dPKq+iKupfWzAyMYMvt28VMBdu1hxWZqkpUX84wmH489yV6MyJu0HalDMU3fCKCFdUDTvGrnng6Zun0R29Zp9mK2L8gNJBM7yEuRr3l4qQaiC6P
YL3vMpjZA/eO2aDmjv68BcvqoWgffjP83juZ7QQep+PZiG3DfHP6zyKWpTCRhfeH99ZU9Id4KkYj+jnRS1WcqXyVrjddaE4jb+Y5QsoSl13iJeFwYPG5qoRDuk3b9BQz
UU/ZDbBAp914Bu5+RtDVbgmbzPExbhQpAgTRi/SqjyArmU1w6HgK9W6S+h+c8ESg2y4yIzJ3z18s5t+c2z6qWtjoO1vOhor4qOg9H51UJSIZA6eS+JAc2jKXJYWHJLap
+mPD85zaqxeQm7Rrsv/Z4YvbiIhZmebL4klxwR2G/j0uhyOrGQtPuxiqUHn9x7ZdEu78Rk5tBt2oyD1BkecX0tH29/usgLAxCOrmGwKrch1hHzh21lGAmW5R6VsUDozw
fI7ORZ64mVVXxkCpST0hp4V4L3RWgmcgo04NcNcO1cvCouTezGUoCLrkUtiKWJwCIz5UyXPmhOz0s67qs7RcZv1SF5sjmE4tyBwHTdqL9CxrYPJD5RGz9O3yjcArqoHi
Z7QqaYv9Ljx0/YEtH1w+RSzUABuTt8JjbK4zMlNz7Bx6vAbZAiZwKMo09dnN6/XLc3OvKwnFzWW8zbxV6ByqrffWVPSHeCpGI/o50UtVnKkpARS5lnuDBiVda1I++D3t
DbiOsiURLiPQ9Ixom59nmiE9m5hWnJ2W0KbOJp4O/kNAEOY24sIkYsZTL8wivJJEZLpolMta2oxNtNIEq43rtrtkNsMyfYJA8h+As2Sioe3972o+/kdgA36cYmyOyGu1
PLWhKrKKJZDmJtPpjyXUk+KMmvcPbVr1uChz/GSj7/Le4totIubw06TyoVSkrCqFj7Ls7HsreVSa5HrOSLzm/qEjtWamsb4HfwA0OQbaDawjoxk4n4lTuIuj7F1RIGUS
ZrfT/dv5ewL8NIG4mrf4o4+y7Ox7K3lUmuR6zki85v6lFAkz4GXWXyle5n24Ydq3/qUOQozTq7BIjSo9+H7/jP3EsPnRStfs33S4TGRDQq+Psuzseyt5VJrkes5IvOb+
V9CS8ecDodymaRtcdHxkn6y7AieKG2XhjDpp8/u2lNdXEFxkBVw1rVFLsKW4yOPEwpQj+G+ZygQ0kT/ezjhAJ0wJ4SSLTnBKKthhuWw3z9domxwyFy+7q1MYCJOSRqPG
vB91eSiC3IatxPCUsTBgrvKDZtNwX4pcjNWRivOJ+8fZ5xi10nS/nBEjGb+IC/40138JmrxVKRKGUH2AsswEumCTL57B0M7fpw5GWhaF7e9v9blmYCDKG13odfWPV8J9
Atf/OKpCfhik6XOA9rm9mj70tPgle7D0F6Sd5GjN2C9jkMyR7aPPIPT/tnC4VjXhI4Rwnndz+8EAZDbRCrRdYu2YKPhJadyRw/cvrEUeGNwUfNHgWr20lx8G2hTKnAB6
xaW4MRaBcQCxZlb7s24W/lKPA7ADDR5EHmJK9WysBvhVVq578Yf5x2cCWAeaMAxlphjcFkOE4dUchY3HSd+Pqdp0XCZGCk/nYDZJFhWuMscHPFvt26rEpj5nFnP99lYQ
pK3V6n+9QXje48ABidFbYRnMUeb3QtjiUAdUSOhcaDR+Y2+MR+RyJFAA+iH6dnpix9SzF0sAoNvzjsSywH6Z2m2Dwo4yUK4fIz77eUqkTawBcVteVejCzt9VjrSBKN6a
RY+NMTZjSHqhQPSD4THWLSo3VkWvkS1wNuDf2bwNcDtgkBNOGeY/rZs57XKQRlrToJVHIi081OPoSNP4bUmyrT7+kE8eLLjdaoEXp8B5g2FQW/HU9vA3wSYVp/3HfBUJ
cxzz9qqPWpPc+ipP1ggH27KFvcRZFwFT1r0ZTbOxH9r7tx3nieDnfd3MMWbqv2vq9zCwBi4J8/tzFJwoCBNGm1O9ZZjQaweM9LnBwC0H8DTk/6IZJdEjefhcHV0jYhYg
O4QD292CrDCnXK1AJKFheAtKOS/NJH9xAneWc+69IP08af7u3aXSEGDj4xIRhqUZHUbdIPN8WbwgW0NgY9avRk81GE1D/7PpIf/Bil3RB8DydWEuLRBmGibOA1GCqdbN
QvQrPx69ghjEfZB6Zb5XtXs+pBRP0tl4j2d1qjSQoMCh0JYK36HU20I2e7Th2ATXE5rHaOCIv+cr9h4f6eOSAmbj/sXSxEVBFy/UFYPfeDCqDNdJcWDKXnyf8VudGaBd
dmMbHdMW/tRki5G3Hpk388oAeLYc0Vdd3B6ySUcN2Q/IWxPKA1Tfj2XNfgebSTUy6kPxGJmsYHFXAKYoUMYJ0+6syo0rS7DScWv8ISa7LuxmTwPWa0AAhbVS2H2s4my3
vC8fVfB3XVPNQQsC/epbkiJtlsZ6L/3TKyn9LKw2YcQ7aDGYtkd2N0gbVo5GvlWUswmzzw71ncJi0KZyRTXHRH7bO6pHllG0lLEVU4amiq5IN2Uz6Pxg2+hgtk5u141s
42tPw7TpaNcws+pNw8tNXzsBXaJz8yADCUoyEJ3nP5RVyCsmd1GmLDOczl3DAnj36Za6cGRAHtfLNE3BJwsmohnMUeb3QtjiUAdUSOhcaDRFkOzrItl/VpZ8mU5s3WZj
lNEHzTQkAG7C/a4MEfiPrrkVWUFpFy1YAGD8sx33AtROAFdA7MKxGZP96qYkR78EqjJqYyDySnealSXY4HKV/ldWs8mgMHO1AEaYGcepNGgoE9Mcz+7SjyKmDpVzIkpv
961Kjjok0iHYUyDIOR1YrlCzlYD1hjbmo4fHvlELrPf0VbYXoBnLwmFVJNc66J+Q4RV5gG0ei3t5gVs7eUGIAVUzScO8+IGkZplG20GhNi0stEW7lPvbPK/Qr5Xej/0W
BUsdlkP5SAKfpZMCzoYQyBy++RIaBweXlub12Lfb8wzmfBq9HJURpuee/joOXJ+2tgS7lVXpG9F8pfSLbLf2u6p+z5zeYG8PUggdue71hBZVyCsmd1GmLDOczl3DAnj3
6Za6cGRAHtfLNE3BJwsmohnMUeb3QtjiUAdUSOhcaDQm4yCoYb6TIFc9X9XvjTZyMXwkzZLme3HqLHiIDbglT4ezLc8yqnBoEZJIZZR68vrQxI/OvcxeazATqf2OaqbT
8yybqd8f9mfsY3cspq1xBGvuQyws0jl0tviKzckM+Zw03CaNFarwGljRlGEZpuEMvqczX1QOfex7XQLn2fiD9Gdtedbq7u7U9PYdzGAlrQCJnOzfua9ILIj5yTIR+Wxa
Ry5BYvxVRYo6pX23Rwgl17aHvpwPxvYoHj+paxvpwPsB3vQnEH+DjFLjVc+FA7DLytQH/K2Y/KzBiOFvCO4AmtdPiiF7BWEzhum9GrrdmrdGbDAq5TQ5/si/JjyPNHPD
Ns+VYRj0vJjm8rcE4ogFB1dWs8mgMHO1AEaYGcepNGjdnFF/pAXdg6FdAIyt1HS9moD6WNPgrEbgeUapJZOHrbZWhWkU7DE/vgKO39lTO6CfMTyIBVWh3AWkcqmzujNk
V1azyaAwc7UARpgZx6k0aN2cUX+kBd2DoV0AjK3UdL0HSYxe2HAkqBqJWK97HU01oumqh6qAJTcghnCy0XUkpsXB+yrBnUiLrfPY3F756Rb9ntDob7I+o1UHLZMPxUMa
fhE0IePkoIhyHfd7sPUY/rCcnIkeQVULKreNp02mpdIVBMwZYgesOnpKgAFx/js0fhE0IePkoIhyHfd7sPUY/rCcnIkeQVULKreNp02mpdLDuOJ7pFvzj2fXn9PXrYcw
fhE0IePkoIhyHfd7sPUY/rCcnIkeQVULKreNp02mpdLK+1pwF8simpd8021tdtshfhE0IePkoIhyHfd7sPUY/mBaw/I6AzK76Z0DaL/wVBrYF+bMflkeO+sJp0dZ1qpM
geUE7x5eBm0ilUw0a1vG2dBiHVtAUGeh6ZoaWAP2gKPqJhUGBQ/wzU8zMWnRvkGTmO44izd6Rg9Q7eRcpz6qAQ73Ehgvxyqki+Z6clHpSRRLd+s+/la7IWn2NsRHiIVl
+THb18WxGS9QnjNz+6Ywp4iZYt3rbWEoV3mtQMQ3ZRHjMxzAxxKdn3aglYGHfxMNHdd1MZWA164UQBUC/B1l9tG77uA5FzeZq1ZnMRm00YxIyeep6O/Mpu0k4er07krL
Uub8Xm7fBzBVdOpibqTuyFCMKw98N115HfFOZXGRJEIc5FqmmgIyXm7o9jAhHVW+imXHwpRak6ScwGsZp4uEuxaZMMdmcIx3umcK8L0g9DZC3n/GHIQdAm4qamRyJRSE
DP1sphVyYv4n95Sk6Yp3OF0tbcTuBa/zIIuZpxNdtzAxqgahb7okJbplKO9Ebcru1QkIlKAFH5gbMl2mGSiI89rK4ZPkdQWKR8Jgr9VPS8P80amlbLrMBbJ3WsNhlcja
7ZAtWbCeVEI6yCqugXP3zfxMVFNIqJMNBec3EFBWe/OZxSiKQmgQLvA7y66kjf3FJG4pyeNwg7b6Dudcnwcd3Ecjhd4F+cs4205jcsRsBCn/ikcxnl8c+G0SIcY2qRnK
sirgwLFESImfphraWkbSpyTLJ6M66ro7uyVt5AadjIWtX3cB4G6JQtOv0g0vD0vS9yk7g/iwMWYQAI+kPOD8mV0tbcTuBa/zIIuZpxNdtzDYIJ51J+qT/Zl4pSSJObEL
7EXOGu/j8vMenfeI3AE0TglwCnwNo6AmtELSgNnTz+bY6DtbzoaK+KjoPR+dVCUi3eLeRAYv72L6/S0/5QYdpzQDONFLyQOJPjWRHdnIh69MQ+9OME4tlx9ra/ST2yWF
Xoa6EVnoQQsSMGzbCjW/fNFo+Fqt+VOnd53RNNQxi2gsRhaNeJyETWq+90VTZWfKlShWgJzQUbnO5j2K35n2mGNQugVlUbamHK75Fmf2qly4YwxhWZg/DfyhIqO0lfu0
hHC6BVXmqgfT10idaKjnO0xJ9OFCAUY7ftAkbwLAl5Ts7ZRJaEJ3xYUV3/RFOiYr9jbz4lAqWhHab8v4YU71kESFKvEZEqqlOq/a0Um/ysDn6QLqrsYS7gcVRMbnwnkp
jyFT+sOBr0i0s2jeauD6uKB2UL2v/j7QJ0hQe447yVWW84r8LC9B4uhQfQLk1F1j/R//LkbUFHm2pfPkwxssLIFnLJYp5xkrX0pJCZ8IxWp1koGYY5Spk08N6GPAOiyE
0+sjI2WVqKHRFDrQkRjFG9TakCv0ZOAwM94ijf1TnYIawo5tLIP2DLVPlEA1h9d1iOuceqxdFZiJ6ud/3e+XFtjoO1vOhor4qOg9H51UJSLd4t5EBi/vYvr9LT/lBh2n
n4Gt8+8X7V2RYSIQ3e2IZ29kWWVzqSyf+I1rPjNbt4r0VbYXoBnLwmFVJNc66J+QiX/GYbYhGJ70Bg7NEON9z4CmNxzirTYd7fXcs4sXVITYfhu97vpUfr2++uJvctK5
kQV4BuJ3Ng6r4ov/SP1XG3W7+kOHYU3+2rmoyqu/CZR6cac5rhmkYj+wAu33UzzjhJLhOOB+JXt+WwM5+3oMm8Vm0pbXmQjWooa5jiuDxD92eJjk9EYN7N06n62i6oDh
99ZU9Id4KkYj+jnRS1WcqU6hNZVjh2rOBKi8mchUALBvO/KIa8XjODTxAftEuN7XU+2JMUrVQLqzP9HYZcZ3AokuVtY4ql2bwagvy7Y1sz8vt0X76QeVHKxlYvhcVgeg
5Fpy8VEMxaAjZwkS4SOZu+dfcFErMw+SYY/pHAOkxLfzj+K8TMdkjDnDU9uCZ1CVUobzOkOH9p5tSStxlKhjgrgHYBeOU8+PB/BZgaeDRgT6w1Y6xLr7stq//XVir3eJ
F61s0/IyTxzh2igsU06SZ/xMVFNIqJMNBec3EFBWe/McrZp7Y9cGBWT1PR5nOiiwLG12e12C40jtPF3eT2Poq5/5JZYlSzIWeUYgMrSqKrT3dls+OIPLxbVlgYGqgwuV
sYwWIk4811cVORPGvRyrmN46TpUSxWiAOOr9vMGrNS9+1Ox8vZtPXSuu1AjTBwlIOH0jUHa6An5YAhxYzH++wRSQsC8Vs0z1i64PpgqTjgaSKSJxOLGN76eIo/MDyErc
Y3pLPGnMEHj8qazZADYd8mv41SFsGPNe8X2SdKqlu/dWO3jLm01wLRmrH+hhVXXLPeoWsGwY8wGmXjNnNNJE/Mc3WHuQ/HDpT+/I+FEGz9XQ87KD7qYVpD8a8dgROe3a
dD46XOsaf67vwBMz0Ua/ZwRsPcUq3nV+saWjN/PZTpdhdqXq2b+AZUCwfXiK7bQbOz4VyjAcg9Zlj+cwFwFDXm+3Z9S81YVleD+90fiLtFPpDwEEZvyPjqh4KSNVbSCo
YYasSZDlQCyhNLHNo+JtCKV2F6DHdvfWswl9yT7MqgI7PhXKMByD1mWP5zAXAUNe6iKDFl1i1GQTHzHVu++jR1gF9GkqvI3T532KH4N1qB2kClKN1FMVnNfxNyF6FNRf
lwGTxSZbB/uvgmakt4kn0dxw11ZoB6xgIa8K+EwUWG+5CcbtYQbBmrjXDifj9ydgQg2OpKTz6PORwdffKfk9VfEN6rRk6nW6KQsrO9tHpR7GEk8FPF0dILb/oBJBXjOL
4xFg9IsPGABCFjL60MwXA7kFNNw0xEq+4jre/PG9io8e2zEgFUiCziWbMENyBkrZnKCekFiJWUxqFRz7Q7nJWYGtQPQJ2wLRTcjuy4umckRgrL3bOrjUJ91cgceBjQiL
OgbxbjnHH1TS2qbUCjkJxQ9xsc/UJNwMWEYrszL0F8/l1YhB4W7gMIslNVqN9TC7OgbxbjnHH1TS2qbUCjkJxSJAT/u5OTFKiKxQOL8MbZQHUOxEX9PHYe7cWVAfM7k3
OgbxbjnHH1TS2qbUCjkJxe5YyD6md3ialdQ9sN/lZuJk58NvRg5mXKM7i7uZVmc2GADDGXUJLeF7BSj1OGNYxZNN33Oj2BdpzaKaV9WGQv3UAY5GIQ/T+PZR9NHlh3T7
LN6rpvei793m0DnDenzA9GTnw29GDmZcozuLu5lWZzbjmcBI541sjxC4IM94QLisS8EgEux70A7NVBs/T4hvzGzhvktZZ7bxRkKNxC7cOmmAUEq1a3VPGPZeROrMhuTy
NTpfnag3BoKoe8AusaIom+wHedLVPHtGD11TbVqbHNzMUMVJnldvRz9YKl+K0QL7ubNY4zn/kprTXnwXk13MNCkINysCNi2aVp7J9/SQ+vxdM/TdwD/TwJXxjVTaFxA9
yBpkQXReIyPI3E3r2faod3EGdxDyxL4mAqzOEoYAcs1dM/TdwD/TwJXxjVTaFxA9PVrBOch3pupRUcm3D4/AeNkUkRhUpu1xxYYmXZZgJO3SEKPHDZOU7Goma6YiclEw
+J9h+KovGBMCYQa/Mj5O9zs6XGoZw/du6EWnUhX+2DQJ7J17qpAxjDIJxLeYg6u7EuIP6HsGJ87b47t4LupJfTbV513lc3/eEEYp5LP+NBG0VJxkdvJLGZ0+lXRPipmV
FI9pbfT4ZSpGVpVtq/2mFgDdEWXiSennOooQrnArRC21Kt3st+raasjh2v1+ysA8x7WCSwjf/PCFkEQS7KxmXoacL5mkCJ5Zc1xiXc2V+A+J7jwDaLNLj8xMBcae4jEg
0TooCBZYm9AePULi8dyT9LTkuiO7vlzj/U7XtuTcpubhuDna+yvzwyzF8o1d+Qx15vqifn1EiiXoX1EWViwY7JDdT2rcUC5+gEQ/BhhH+/V2MMc6ofMJnaq/uazEhmpe
yogm0Sa9h4GMq195YwJtiHUN0P6/yW9boRnJipB/n4mOq9kX/mCNE0M04qkOo7NSJnuQXGnFuDT5U89ZCHwHOqn+t15L9rtVAGdJpQ6Pypii/uNg5LVUb3jDP5/ozVU6
l46UbFUEThb4R4I453BWxqL+42DktVRveMM/n+jNVTrwDpw51liYfhRqM+Xm7UIrov7jYOS1VG94wz+f6M1VOipkwqz8X6utn7tva+LP5eNRxZ/iDKJeIXyl9Ihtj2tm
9t6tKJSvPhykNwuwlJHy01xU2AfTmqo1wI54SDhtOe+1g9IzQ4DM21X8z6drZUCgupScgm2uHxKCsC14NXilhJZ26fL2w7VhRUm1wtHHZQnjXEeJ596f+lT55c8ZsKFE
u0buPNBFiSgZWoD5SvJKFgF6SW4RUPAEUN+DgGBxeTwhrvcTsuiW3HW4BL3HspJGIuwDE37aKmeRwaCE8aLesoBdUO+RlJE6THC5cy1uALkNfK2I67sFub68fGxAl76C
QnBuiA3CRhD09r6nrhQc5CxdXhagTaIacxM4sr4xcCTUNMXDjjkuiraRYNBsUm00nqfcwrqoZa1F4McfK6BTNMPsb23bo6xdQchKw/evsqcfS8u9DiOC8ZfsKVCD+85B
lCMQqxf32re+xkXdGL0s7f5FoV1cfN+elma5lGb5dpqG0dNkJ9+BXaYjA1zLc0N1r2QUWecyZbt4PCAKy6dyN0g3ZTPo/GDb6GC2Tm7XjWyUexs0nwUFls8gEcnYS867
WUnuNYO06fkSfNyw3O6woi5MUAk1kBtG/WOIbORF5RvkxWl6rZrY/wCJhm6JXEGqgMYX/FpX+4MpfQD7eXLO+Zau21EQX7GYn1vIorqIUuBmcaBSQeqzxsd9gJ1AvidD
vy2Co3eqJPKsOleUQuk86vkb5RvtYRjD0/2f+z6HH/Mpl9EP9mbQw3RNcnVs1sgNd2/+109pxwxzqeEjWhHDRQuPc02Yji5bgV9311H9OkC2ybiFQYBtd5rFY7Bz32OX
ycKxCSaljtyrJQ0m3RwZIc/DA/UCc+zVaTCV7l65mGFVtRmRefXC9lsLr/V3lflO0TooCBZYm9AePULi8dyT9FZmGdFV6HzK3UaIskuRvxksPv36ao9XxNo/raFihewa
fMRs/8BOg+UBf6MAzWk1y07Tgeocg5Q+SVhPd9oHvqnZHXgiT/T0+p9ZnSlLpqnF4xFg9IsPGABCFjL60MwXA2GBvykcOP5DwFOG5+0By+BCgWN/UWQ3HTRXF35HDqnk
A1IGUgceg6XkmkkB51nUzjLz7ahn6DqkUEOU+18sFqh+iW9oMCFOGpLWb9kyOmMU4xFg9IsPGABCFjL60MwXA+AwatBIAJrS5NlNJTyoqTdCgWN/UWQ3HTRXF35HDqnk
u1lW9TZh5LtHC1DuTsMS1ZT3WjjR1oaMfSycLuRPtcCnxV02cL4fR1UkkStbVpgM0TooCBZYm9AePULi8dyT9FYp+J49YJqw+GWZzq+aceAsPv36ao9XxNo/raFihewa
cR9rW77AII+nH0nSdHYgo/yyH2vvb1WFwg7t0VvmKdCil80oAJOmYjRSWP74/ZxQFvkSEqv6hhr55m/7w0G0DjTj8YdLCA65XTN3rhExStTySzaaTSRKd9/aaZL8WyU9
RyCpPeP5uYdd7FkxuxMDa0TDYNlpKKOMXvYX90KuaNqUVAg7idpgIf73Swca1V/r9I5oWlfIHcPdJ2IpTHNchC5fmX0HlZVhJc/Sx5TQXrvr7Awd7XAgQkQfQ7OnLuMR
/sOuFHGfJ+11twL1vaOUESMp0CbGh7iLy2UP4ZKVJoLBriAAcDUKVCenkL6hb2bODDQYsF5rFiYmTstPpGTgwGUvXig1hiXyhDj94sIVZvhlWqhg38YOk00uC/qSyDHI
aCwc2uZjuIS3Q8iWqdaKTNq1ZKLMpFAvPnPRupyJoyumy0u4bOxPJkCRw9aEAAfQAYl6PIYb4dxJl1OjfP27St4V6m0BRJ21FwQXRo3gMbJ3lBHJ7k0LtnIMRsNjdKOq
tMcoeUjNre+vbZLHpI4vFlnFBLeRQtZbIeCwOSOPyV6UcESzfzVChPN3eNfRQp18qzojJHxV7MjtcCiHasvi8a/cdO2byJ8qpvYfxo6l4V/cNen1K/+PhpzjsLykn8Lz
PHPZuTupzIZ+IJW0nEo7pYQ+ac2JI1VCjd/9nEcZJgRbZkMDSXZhcRvtJt5vPBKsQbMzfSx66qPe+BZa6gf/Tel2AsEQ9kzeLUbm1VyU/VK6MqrstvmLGHlwb4q2xjYL
WRHGqr+09lgDKWhj5yNqmwKmx474stB+aY74dRgKOnW5FoXYF0WGjjFcB8eI5KlK5MVpeq2a2P8AiYZuiVxBqrwW0GDX5XBpimLBTfVBGfRZpx+ugWeLYAFLc0ThJ3BG
YF4kMUrq3SSzJvlQXaXp+NrGJdq2g35LSODANsztn82psymwChi7rENQpnL3eVYCa7iadA2o9BJ1n4EB03razJ8FmiTCF90lCl9I+aAv4YEzQUu+El2b4wLNZl558jWT
5YulsJuxllqZGn0v6sEgA7RUnGR28ksZnT6VdE+KmZVLfgXFXilvmwccp2RGqYAFPAN/PNCgmIrf96HNaRInnW1NJyull9bUlPVR1ueAUWmWnTJr/9PfS2jsaIIAZ93V
VfTzGeE6sjM6aEEWhcTrgwFeBog9tG9Hg70d094l4/8zQUu+El2b4wLNZl558jWT5YulsJuxllqZGn0v6sEgA5ygnpBYiVlMahUc+0O5yVkr0mTaNQ1FPxdNsV0Hwkl9
q0GrhY7xoOWuy34hjdC7H8mRPHfzMmq4uJ5FmJSUg2GroKIRXaJXa4xJBtiO9Z8zPvscma9cfn+2u4Lf8mRnoIA6PllG7pC6+KpWpWFJWSzROigIFlib0B49QuLx3JP0
tOS6I7u+XOP9Tte25Nym5nncEOIjNGKJYSCfCZoH9IAO3+nYmei3D6286yNXY+E93Hao0d+w2I1IGlk8Qo6Q0umm/bq/yLMTxwSVvN591Ebm35guRwVJZxAeqkoB0wBH
e8teC1BfQGUeimUV0/ASBWuOQEBPgr0W7RC39cz56aIE7L+9iRSyIwt6H6KWop4tGuBgOQkCBe3hxCWTX9qVbc24/TPjxyKqU43gGZYe0ScO+AK2d7AdoFlPZJ1WM/fN
DaCxRn5y2rEHEv9pMyZqi1PPSxBcfcxVu1XdxnPQeUps2MNFy/ATUGga8+fIVGPY+YkE8Vpv2zFOdUlHXG1767lihgNtTaXYgjI1KlU+6LIybaDR38O6jBbNd90LZdbz
2xDCzfjQZp4kwAcvN9bD9WHU+mLMgcK9sHfDr3VqGI/+WNCKwabbQzJjx+iJHz5oUQBGXQgZOpOJVE9bMGqbO7VZcX7l6yFrhCIP0O3ArML31lT0h3gqRiP6OdFLVZyp
BvJdWrSxDRR+mW3y/C1/c7/ndwKYjnFyMreRiLYsnBW5YoYDbU2l2IIyNSpVPuiyjFUYIbTrtvL9h+HTQcHFhAA8zi0SMruJiw3m4wuAjfyxTF6ESExL8sYsK0I38pXt
lxhBREdPTS6LNg7VeEK1pFgF9GkqvI3T532KH4N1qB2vRCaMKfb8q26yR6NXzAUfc9UPBNdVnZbF8BPlF5coVF0o7A7sb73S4MrpvKTXXE/SC77SyJmCm6nUDYygl8Fl
y7pul/SSjKkSFppMpArJnFHHNxHZiXu8SV5haz/hwFI5Cf7PbuxpOx/n+8EYnKzG5R44Xz+rTyd0vxtqRPBZkZNN33Oj2BdpzaKaV9WGQv18hz4sViIAFjhlAXnPznmY
BeKy6yRYiqOWkZKfpthNjVDhScGQMisBMGbux7SOpXx552et238vJqaJkbGMsJgFAw/iX4OpG4kn50NeuhPHZ4BSodBNruHbUYfqWfkt3t77Ls+V0AY/1Sbs08TkiJYW
TyJQMoabyTaGZ/Hc34y978SYE9KTQoJnkpNUEuMBl4HY5AUmaL5akcS8klgJdJkLkInkkT5g8XTbEfUts25QKpW4QpkZi4BHbEQbvcC3hN/dn61KE6lRri0QqaV6/H+8
1tPwbh0rHsqX28rLT+OtJz3aX64gXpzElitXxoWGK8y3ocA33Gpb+4w1/jx/e2VARy5BYvxVRYo6pX23Rwgl1+5YyD6md3ialdQ9sN/lZuIh3NQQuvo4Y3wIDm8OMVhR
26jbKj/5pfy2wm+asRE+AVEzZMDP2P9u5V8bdiKt94odDzvCjNT77i2NpjkAPOm8pEKPbtJhoYNtE/Mv99bOypBU14sK81Vyz54tGhCAuDzNzqr26LBZADP7KUNUK0Wy
ZY8k+mCwegsW6mqrOuybz+KeF0NkCKzNLiDEVw/RxNj1Nb3bUYVS/Ldo4VGlxN/2yZE8d/Myari4nkWYlJSDYZT+kG+uz8Y+khaLMd+ejR6R04bieSrAPaHaoFSDskl7
7xNsfSnawPp0418jdqIPWF8S949U5Mr33XZDTu7g9Z3dN/87QUDHUQ4uYgRJkyDdCYw6RehikSpWMnUeb5/v4HUGRs5Z6q78pGkU/Me0oifPZXmZI3y9Ry1uHrwcfcSs
9TW921GFUvy3aOFRpcTf9uKMmvcPbVr1uChz/GSj7/Lww/YE/oTw+Jc3rIDXU2624Sfxrac6YRBBS8u/9JwWfe8TbH0p2sD6dONfI3aiD1hs1PJCF1naFak7R35td5gP
HFnRz2MQdfLjJI9RJoIdhZjQ0tiuNAp9szp9dU/l8SVyh6I4fBQ56vTtM00C2UmzAfgXE6TE/9kD9bzMz6A9tnTkBpTX52Q/OHkwyWCxAIpXE3UUzBFTw/0Ehr9cC55d
dJuBBBvZlSde3VhOTgDmf0EZNVF2zpVXFHcYzkKIaFoaHJ5097bomfKPFSwaVEYElSXZ8lPw63vBEw3Zv4b/myGPTUuZgaW62cwg4X2SpLSPku3lBRd92YBUx9asJzV0
iydldj7wohBhDviqq1KbUDkL0CWwAc18AUbAjB5d/fPbEMLN+NBmniTABy831sP1zva8SjMdbsowSwakNinq+iHiIPGGXZ0wMXj8mh67v83ccNdWaAesYCGvCvhMFFhv
IjE1GaB+QnvN5t/w7sK8yvxe3ys/Z7A0Akzc0zSOQD9Gw7NaCVZxuakZYKCdm29WtGod240Fg0uv+Obc5Xqew1L1bVEYSLCZ0J/fAabV6Bwj+Oiii3Ru+r5VVAzj0K4g
Ln2d2Ok9xoyrq4KhlSBP0u7U7X+BN0djsxRx8VR3xBHdnFF/pAXdg6FdAIyt1HS9WAX0aSq8jdPnfYofg3WoHRVC632IYayIYTEgxKTAJKkucK6IgPfEkwHqN2QMFuDI
5XfN42XVmXs04BAlOB50AUAyFOnSfcqe6PPzdyRxrhTe2DfolkiNM3wPtVD1H9WyLHI6DQTLtQi7aiPKhw8s+VhKkSbCB/SjAls3oTX+D/vnXkNVtW0xO65Xi/vivL6Q
We4rnPPgwS5HwWU4y/ZyC7zzFNXl2kfLvtbc6On/mIUdveyd7tK5nKILXXmTISqhaPSKt9oY/jq/F8AE2WL1fwQgB1UMUahCNKAq62KTL520NpbYKr5fovvwdq6onZF1
BCfiXQSQK65L6pfIBBsAISewlS2VnEIr/IWrW0pJ2dJiRBcsgg6zbOBq9EbneWBvi5IpdFCcD+FVTbzsNb9+2am5WefJaGa7Bb/rR0CQAFmrJ4EQs4g3bjObo97mueCt
l7Gz03C6r9t0weyQ1ZIz7YxkX/PBSVBmP+9MVBUCSBk94EIKK9zGm8DFmITLeTHWJbXiSwZKGCYdaEKkwihGbFJG3c7TY4cr30VCNE4mV6JHCi1QFUxtj+gbgkEOrQJ9
EOt2SXQT7Im1yPdbr83kBMTmwmx5Q7WifocwqIsXXCMah7NF3mX1cmxNBYDluMCz5bvLF20j+fvFU4n6Q780tZDdT2rcUC5+gEQ/BhhH+/UR6Zbk7p6EsALLBNO/hdoP
AieWUND8t41BAL1b1Ktw5cJpZQMuUrlca1Zjc1jgm3YsKdbK2AM8Fm6Q0Cug+hnNR2xPEdIx7xRpEQD2z8jxgVVk6wxY8O8dK3ODSO3H/6wqFyA6BlBqSq5yqXx5lsl9
KJ4lu65F8j/1yMp2iPJBPVPat51hnt/gVLpOqme2HYYVEoyf1UwJIJo+p7QJVMmGbpnunq0lpLRBRgmwE+GSQALK05kJnk3i4d6W3H8gEFGpe5Miocy10XwJPX+2Cn2D
n5eZrY/05yVhJUloM2l5N1K8df5rFex8guT0Ahu3IJz3HL6Hjm1gNBY2Q7JGt5y19Y2t6kBXU+emBjFfjiVPhJW67SjI0hPdhnwl14n22h8MrlPLg6VrhQoqxHHU5vIl
2kaPBHp457UQ/nN7TNsCyNFY2BNeShvFWIV9UzEuh/4biJ/rRqeuM7LstK2S4OP7MisSpv16sH3gwo8vXWPV1JRCskm+rDpugcEXoM4YK4miZvl29v6Cn26qOUx6JyV5
g/vcFZLI02Y94vkGISIdcl6LPD9jk/iKr1mn3ngJj7ebQoXuGBOyndVud3OlmA7GrTcW1k1r3OAZIIBnuJI3zP3vaj7+R2ADfpxibI7Ia7VpBE+a6eI40QGJzF4XbQ3n
VlgSHerAtjOa0luIVs0k/6fNCHpNvD/m7khP9YRRpXerRCTDwMXJ629SvvpUSKg6ipLqqR4uf+qQcmsdZMGdgZjQ0tiuNAp9szp9dU/l8SWjT2nHMbjesu0AekuRxaxQ
ijKijg89e9TR2vAPcYPIqrsOYme3hxUcR2IUjqsI//BIHqOfEHsLTpHSbi5HZyKypRQJM+Bl1l8pXuZ9uGHat/6lDkKM06uwSI0qPfh+/4z9xLD50UrX7N90uExkQ0Kv
csBpDpAp/B3B4Lo7qJyPmOPe19PM6JAKS04VV23BZi8WXqJLZqev+Jt7275yFil9Voc7X3iB/jHtnmFVfzgXFhgAIbjNjYvaH8g302shjy5ntCppi/0uPHT9gS0fXD5F
hxJt3tOwZHUnjDCDavcGwxga4qWAUYaQ6Mj9nhKDYBmlT2Mbaz5BAbqTS0z4aLSnCYw6RehikSpWMnUeb5/v4LJj1qD+oo8M/c6p/tywHi0MYaNhJf+YmFRl0wU/BmPW
lxeMavO6RVGnvlnlAiVMH6pmB/VKu7S+Ay0kh6oSkxsXm37Zoabts+RcgYi39T4HXIxE58QaAWC4TGe7YPZh/VqBII5TSB3KnkuVdcKkzgdIHqOfEHsLTpHSbi5HZyKy
5Yvc6OYbAmNslj+iZuay8AV0Pj1N1eAO1DIVqnrm2zpStwSYKVk/24b6qxVbFnabaefYish0it8sn18CzcKuUshSnjKuyuSMkrh/00ZJdZtFFYM0p3YH0lZ7bpzWjUU7
S22E4gg7fIlH6gNoFoJ0Mmr4GfI50BxwEl0ZYIbJgUZa8bCulpWx3eVkwqmOM70mXPOyDk3IC0mk6GbfpWB41EfUM9h6hf9RX2wpjGU+SfX/UfujnpxdAWHx0K/hFZPe
iDU+YvQmB9KOBhMSXCz0G6Qtlgvq5Hp/YwOX8NE5+nkAcmBid61FsUikVpKpE1waMM06zAsD2tJ1Gn4dkASwNvmB4B72BPePxSsEENpraUzSQ8lNBsbBYtsgVFDpZsLg
mNDS2K40Cn2zOn11T+XxJX7SbGijwGqL2sXrrgJEvflVE9SxMAoRi/horv7DbpJrpAUejK26rInmFr4gzopwi9uo2yo/+aX8tsJvmrERPgFTYyTerXB0su1jYcSlJ9gi
dkylbxhiFgitz4W/ouoQNMMBUSLi3Sc6sR7Ti6N7EWe8KrU5au8kYFEBP5GN92N1Ns+VYRj0vJjm8rcE4ogFBzetLlRDfwNp5g28NhLfgnxCBJvWGvk7CU1dslJnb8+i
R9Qz2HqF/1FfbCmMZT5J9SvBj/hOA5h/lb4YSn1omWXsIfBGUt16/CmJfoDwbEiPBp6n/WvKF0PK9Iga995+m8oY869erfmKr8QQyFT4reGt63kTaBmVOQlz8tDlKZqE
lkw2dMNX6g0lTTepn6r6bZ/5JZYlSzIWeUYgMrSqKrSLlHv08HjTHtwM4kOm5OW9PYDI9KAypbc3UJnP9ZK1Qdv2yrZbIQCHY3y8nboRbUZ05AaU1+dkPzh5MMlgsQCK
luO57lvHObJ5/f6l2+2GHzOUK96rS8xB48ZjyRZy2f/jnJULoIe9RJ+p7mWVd/U8pC2WC+rken9jA5fw0Tn6eQByYGJ3rUWxSKRWkqkTXBowzTrMCwPa0nUafh2QBLA2
+YHgHvYE94/FKwQQ2mtpTNJDyU0GxsFi2yBUUOlmwuCY0NLYrjQKfbM6fXVP5fElgPc0Ulpe4V4rGth70LwoQZPpin3Z/kLRMC1HGvPWKVmUZsjjgCbqdyb6q6ubQPK4
gaZY+wTWLv2Va5rDtXmPoCEtpyJzxUvTubbO+dNMWvre//1vZC+6blxD4ocDoL2YZQYblsgmDbzJU79AX2xpJQ7f6diZ6LcPrbzrI1dj4T0OsbRdQJu3yetNisJ/ENRb
1U1l8TMeFMz+87twUhG+VGGrlsXGcZ/MwpRiKH/GlXvbmNjAg1IYfBpCGrbKiFQkC45SxKqy2HEkgFef8cgNfo/gV0qLTKbeVHaM2xryM92jI6li53XdjbsgT2kH9zVE
3ZxRf6QF3YOhXQCMrdR0vQYRkjsW/CrarT8dXdAK6P9175fl+ENNDwMHRnkZKtZ3nwWaJMIX3SUKX0j5oC/hgXTkBpTX52Q/OHkwyWCxAIrSvukE0X1IU/ipD2KAEu04
KeTfmmlJfMu9W4YD9bRL9XFTQ0gcvXqvk1d7T2wkurc1gDZqIq03Q2li4N3ttdaioyOpYud13Y27IE9pB/c1RN2cUX+kBd2DoV0AjK3UdL3sMEby1vqiNUoYCVNUFpLg
D/rVVTP81r4ouZR3yRPV0JWlUrHciYtell3CmWzYIndsXu6ZenGomReKxh8vChIhaZ4QC+zsZV310EgP3XEIN0J5XJ2zurzIixuG/mLVRnBWhztfeIH+Me2eYVV/OBcW
U89LEFx9zFW7Vd3Gc9B5SmtALo42jp6Nk4/ydwChsNo7vo7C1WEyWXv3vtabEnyQKnXsiH/cBGDtYXg/+Ds7waoDYQfSNCoezvqr8bPqtkbSQ8lNBsbBYtsgVFDpZsLg
qQNZ1U/+TLtpQRQHXuDh62BjzjjelnVFClGUZeX1nkySc5NeeBWzLXPqBBgH3IdfjgvPAAWX/VM0ZZ2lG3R1F0Ghy7SaVHR8J1uirClsWFJlQng6UkKpYGUam8ehi2/6
26jbKj/5pfy2wm+asRE+AX34O1tNsY45hAzq4LIbQn+KRtkAEMylUJcwo7huOjRuZoL/Wbhd8jLe6Xt7vNvHCMVL7U3bKPDkqIKRV0Wn/vkGnqf9a8oXQ8r0iBr33n6b
oyOpYud13Y27IE9pB/c1RLntkmVZ8vVrxtvAmSa3R0WtbZo2wqLfdJW8F7W7L3iDxcH7KsGdSIut89jcXvnpFs0tWuONOKZGTPPdpRHyekpU5413y/aJ/E/hVXOi4SCB
K7CywJoCFMDuOe94mE01CmEW8yNkAhhGNQ/qptpaKgkZ0pr93MTKG3VVGsMV0Xo8be4K8eN451NU/m/gCn/VFbpAcjY4NNAZY2cEtgbOwtusW9NDtQ2y7rFlcdkgPLET
tIS9Zwwo2Fcs136hmXykRPDJkwYq8v37bjcG7XMu4JUBpCwLDJGSogfZHwpasq/7kP2Bg6tjhRPDmKTS1tSsnGRJJY4rk7InR/dwo4V7KRCpvr2vQM8EkpWyXS3LKuv2
S+C9jwR31B4EFxxXq0GNjBfDLWnfRQJgQ1rw9iXU0f/kpVdz/Ck7J6WDrBsWrf12SwYxj5V7yuLrRTG5qJrv2oCmNxzirTYd7fXcs4sXVITkkR2fh7tsFEruRd7sriOG
10+KIXsFYTOG6b0aut2atwUxxYtpR0JpBcxG+3yMtMTH7cWWtjqjHC2Y0vTybTd7F8Mtad9FAmBDWvD2JdTR/2UvXig1hiXyhDj94sIVZvg5Qv9fcfcJaJzYNlDIiVHF
qZHuNmvGrw2vK/JCmDmLvc9M7R1RCoWsnUI7JhjCAPAeJ5WzZD2GEpiblnhPS4ZIfhE0IePkoIhyHfd7sPUY/saigNYdL3EeOzLxLhxT9yyiX1vgGnK+6RkNEDk7n1cr
2H0MSaZ/xLBaCHRkHT6AsPXKUcBr3M1BDnhoyplDtN7b5TalzmiyWmE+Y6eMsGagc60QRzEngM2cW8MYMP4b7TDWTaUyAvX+UdtO+yuW/LNf0JA1ypW4RKCIrdTCYr66
G1onilvQ+pP6yVuSGzG44m6j49XNuV5YFNcFC6F7MwNLF76zhSFfgexnZhsRZDF2U9IkDqnzU3Au+xtSXEy79OtBWC3zCoPGuNh9++4WyuAlALfx/UklBgBv0bODmdcw
+3JzUImCOQjcYyl+Jk81LCu+svT3JQK3POD2M+Sedufj5Z+2dc97oLtryJKRPWF3MGDjK2e2OVpmA+u6Ew9u4R2juAUPejH1g9pQKSoEHxOFwgqzMhpQJzyppk6muM4m
FY6BvdsZlEZx8vuyS2CxV3Alr3UyX7c04S3KHMHQiryJlIi+qgg8ifhsC5wckVQrY1C6BWVRtqYcrvkWZ/aqXLhjDGFZmD8N/KEio7SV+7SEcLoFVeaqB9PXSJ1oqOc7
UdSut+diUOQapzk9BROlw/gWJAKS/mllbwLodHnJgHQZV5VLJ9YgUbv3j24f4193Xqh4rCYqHXQ93pYeVc/6IAXTAqt7gplayOvqG3FbFWjk+nMdBKzX4TOzmcwnS4/V
GIUhVE6WJBvqnzD//T+M/k4PI1uWyBnZC51KP4wqZWa/QPSgLny31/1a8W7xgCSLtsKFY3PHXNY0RfoK2+OXkxKEsqdER8f8SNiWvYS+AS29dbsC/K6BErp2ps0iSGip
BSNcUxLMoqYL8I5CDgYymsMBUSLi3Sc6sR7Ti6N7EWf4J+hXBHE7Yi47bIIIoShodS66CyntaIqrXwsc1PBPNTKAOhgWgPbkARv2brATO4pxZDUR7gdgv3Qb2i0h82AI
QK6aUMtZYMVCqfRetCxL0UAQ5jbiwiRixlMvzCK8kkTjwRPz7ZViWQacLX+OxS9TdGe0WCJu75ToHEQ221WGJ+dfcFErMw+SYY/pHAOkxLfzj+K8TMdkjDnDU9uCZ1CV
Xc/P0z1IdtHGAruqaOqhCoZeIvFh5t3R5AvSacs3WDPD0glWUpdkuJEuEthFMcCr6Ibk3C1pj2w5K6vlXvIWjebv645Uy/3s9tCcy3EIJrQCq3TOZyyK52XvsqVGbTIX
U2f47eK3vO7pAXcHgdiG6NkUkRhUpu1xxYYmXZZgJO0qvyi7JE/ACnuqFsDsfZQeKbVwFv7lmIE483NxjEeS0Vzu4R55P3bgtmlTrXX1noa2YGUIPAj3YUTGRUOUqTTS
WAX0aSq8jdPnfYofg3WoHSOoV01L7+igawnbk4+zTYakzGOVJDNw340r1fXN/Kzs0t/cDwMUwJChx+VfwTfoHyq/KLskT8AKe6oWwOx9lB4wNIPSfpGUy1T1JaUzhob6
m9gTYeeU0JPm/IMCBezRafSaL6BkeRl2jd9XwA3M4Y9CDY6kpPPo85HB198p+T1V8Q3qtGTqdbopCys720elHhrNYfESH/Cif2qYPexlAXUMYaNhJf+YmFRl0wU/BmPW
QJyx5sKSfmOJKI4bRy9xlXcr0XC6wFHpGpsvYJDSxPEqvyi7JE/ACnuqFsDsfZQe6OTVdnE2FyDiiztZEhE9upvYE2HnlNCT5vyDAgXs0Wmlgd/ns1d6GvIejMzwtSOe
0UuhlA3PO/Njca/ahiW5FYo3ZWm8yuDEYCDdNN+a+wVrvmfC0bStZKXmrVGhpYpY99ZU9Id4KkYj+jnRS1WcqVB9Z+r6MNHopPbDjdRcf/pnHvQ8Z0kVhplr4fnbawSM
M5Qr3qtLzEHjxmPJFnLZ//VGSS72NNeWLSqIPBvh4T5vZz8WHCAWbvpxrKsuEkA/pHLuryMXFE/PRMjP2IrYZ3hCE9Zy7kzJmZxfRn481SMuYpGIjaUi7tf3s84xauPr
uIuX+vf+DrgZVtYnmY+aCcBHGkdCpBEVFc+Y9V217TyQl7R1G73J1Kx0A556GbKOwtWOBlcyny3EL/JwXc3KJqiUZUq0r/px5W+qQYIyYFXp614+Q0J+udajGhV0P/ux
ZEkljiuTsidH93CjhXspEBCJLOS+HkbD+vejgUAUYcESJHaANvR3/LgKNPs9OH+Ktz0+H6Kata5ZKVpZsETs8Dge9io+2wVZSwZj607GOrYGHU8gh+Jkdb78oFLSoqWZ
2Z4h3MDRCDEjtBXMW2w3cExiSNMQl2C7y7UnNBJ54QjCuFEl690/B3jzSHMHm4NBkJ/tv+X3uzyTCb1W+VK8kV2csCtkF3f1P4HGRkrWlWzEmBPSk0KCZ5KTVBLjAZeB
PpyHT3Fs4aOqKV7GAUct2zdBj5lmpcE541vJK2D7dFM57qRqmhxNdfnLS+SNexByidKTNC12B/HZ2wVpJUGu929nPxYcIBZu+nGsqy4SQD9Eofm+0gbeG5popTOcUVD1
+Z8QgjRYOoCowgj/dtNcyHyHPixWIgAWOGUBec/OeZiLPBJiAPn6I8D6J1WjNz5MZOfDb0YOZlyjO4u7mVZnNuUcAJ67m8TFlCa/vVAWkAUBkmwvdVSu/Ft7FGdCD7CN
glekYmtTVlj63rnvhE9pLRe84hQta3yui19rqgzVCW2Fvs0FQwkCPlaeS9RVxS49JXZVEpvp1qFFx3upXUPaNlBPVeKeDxANZj2j6qnbEQZ8hz4sViIAFjhlAXnPznmY
gK50zAXyQN5Xf4i0S/r0FpvYE2HnlNCT5vyDAgXs0WkxwNytL+sYSrTWCKnZibFWvWRUKqVhFhkLTv/mXkgUTitFA9X1IU248F86qtWRXeYpq7c9DrjNbfsn1mofbMFQ
yogm0Sa9h4GMq195YwJtiJTQHhPvwNayxlpz4HBGRkqgahgW6KMfx7j+bOw8U+ORG/QsY8LGI6kFo7BZTfIBzVGi8K+QXQ+b0ucrpT9/ntMfUATscFng9Mdf0aKp8rnR
gAdXtwqDtrkMcTULh34OFPXTmdKhn9z2oWQSwRFXxq0wdBp4CjpOBi8DMTOC0oKQknVfFikngIHMkgsguEwexxb8dZiIRoA4FsHIzIz0y2KXAZPFJlsH+6+CZqS3iSfR
JyE2zgGQ3SNZL/X7OF8oPEKROt3laPXhLEIEG1szlFrXUx1VeVkKrYiVO2EpfJaxPDTdufnexJtddnwY7PK8yb12F2XgcqQmqx35ILSO6NqiHDNDkDk0zU3aXcQFQyNO
7ORcpeBg8S1cFvBHZsohnJk4w6fknIt63IREKmAVaoH7K8tIN5XN0J/mIoGJeHA8M2ELxgdzIXgPRr2al2CgaFbjsPeUkDv9UO3yj2H0C5xlc6Z3twiGxsu9zhYAEJL2
YswXAGLSPoa1xmiwYefboULZJnxFLR+05+2wLmZ9l/vL39CSSYLTvV1DxtvASvtTcsPrXEe/599E1lDF9fAeM0ljJIlaWr6pdZklHw/CpvQfUATscFng9Mdf0aKp8rnR
YL3vMpjZA/eO2aDmjv68BVdZjxqSL151CGwgtEE3QaDZo9WfD8Dbu7hhWC0b33w66t80jPD0IgjPf2SjyM6sB97YN+iWSI0zfA+1UPUf1bJCKZf62Y6EUNqiraIjyuGA
6+2BhyKwcO/WVVzDH3PYz07hgWG8BwB755noMr6iotfF6eajZbkhA+rKmT71rSlTT4o+ycFjNLai+e5fFZWDz15lHBsbx9tqUMG2pvKYLpmHXz+tl75coxOX4KTxKV0H
AN0RZeJJ6ec6ihCucCtELeOJFoBxk4CwQIL1JggAYf3kpVdz/Ck7J6WDrBsWrf12jnv1eBojtsvOm38g6CRlDxJhPF8T4GxbF1tuMcfAcz++vk9xcV22xpv9NWQX4yYG
DyZ/ehca+67e2ay3GyhP0dv8COffLWrpeTlx4oNIFTRIQ1gknJLzv8QPdAIKCiX21SmWPAZ1uv83Hrt8Hbv1LpKEUQ+6bk1aOkKCpoOqwAHV4++M77VdgSMMk0uc03s7
2aPVnw/A27u4YVgtG998OtGYpUNyVSFJdb6NYMNv+MjtyUsOJD3CS85a7SzIsCE7TuGBYbwHAHvnmegyvqKi13K6rmFS+Psumwyy3ucACsi254NMbTZ5Xf3UhC45u4+p
jUJPYuoZ4lAH6xnK/EIFVPPLXzxm+3CRPyg62bgNcaBfT7EYuswDd7JAen+qu+rrVBd5X46AmC9rD/uilGHs3QxTWMgzrVOUD1RG5QSvmt8nO+ol74WXX/rqR6ZONx2i
uaaw7TFYYh3yRC3KHC+WneGCyJRX1qy4yLommnE84cj3bq+HckbjG6ioicZ6zMLWwwFRIuLdJzqxHtOLo3sRZ4vKvqUAxMn1Yx/4GLU9PJWDqcGDNtJN88Ddj8nnbWWj
WqF2uYFqxnb0npWrsAs+aMZxI7T6Zd/jXgmDINcp8DVnHvQ8Z0kVhplr4fnbawSM59vwV+7Hww55U4R55un+v1KGnMdSLU8+0ZR+Cai7k3eyW/nZJ4UDM+UzOn5pnMvC
jUJPYuoZ4lAH6xnK/EIFVPPLXzxm+3CRPyg62bgNcaAtbnfbzS6oySdwHNa00R0UnmFo83c8IazQxWNbcd6dvOfb8Ffux8MOeVOEeebp/r8aEqmnEIkO4cBotuVx6LAM
Opeok1I1+qBzUkkSmfKCLF+gTO1ACY0moTWvgGBZHs+DofiLiNcjDe3vzHcDd8I8X7+AhX8B5vtBzBwF/6VtPkv8RXP8kIjQROwh3OrozCJCkTrd5Wj14SxCBBtbM5Ra
uT68zuTB4b+8oeJFPtzjoSa1IBZPw3oRawcliNfJ9hCufvzBkcpUiwJLhTNlwwBn9C9/1oKEWG+8yEagK6/RbHK6rmFS+Psumwyy3ucACsgGdgwia9kHjjmNOPcQDz4C
44FI0w2yq6YYBW45G267+UphvjfCHwWr+iR5EqPKDLByuq5hUvj7LpsMst7nAArIBnYMImvZB445jTj3EA8+AsTA19evLfMVx/AeRy6Lh9+zFrDRp6AIcYzBhYasdZfl
hg7S4bGXAalLRgixkpf361+tBkWkZUWb+wVPpP0gNCgo4BMBS1zRlrmw0MbCS1qMz53xuaK8IiezCwcLkEjeI9BoUkRKuUJtJUh2HUZH1aQICG2ixdMpDVGJmJfYGfwR
uKppEgO64QpVx1Kbbbif6Y/t1w4PO+QsnSYyzR+OgRZt8fDRd4+3D8j/TuNxLmesN2ZX9HKVDarQaEIX6QugR2DD66azlZu0XneW3fqCOYJFyhjstCIqgDzZsNdD1fuv
gqVDjU1zMxZsSNZW0C6sRCSRcANvA/w/d+13uhe7Sx59PuMP31PIa0TIt6tQS8t5qfJHjThcDYKm5lybTNYEhG33DQj/lNbSEE6wiI4czO2qjEqfOBRVhHIwqZpUm3Cf
AMFSnZ1++bdZ/SH6tncF7/fWVPSHeCpGI/o50UtVnKnlE6F9Jc0Uebz5scHtRF1NYTi08ijj7vm+C3e2NrZUw32WHAJpYtsb19lw1oo+aGhKARC5IE2EUykJY0YlHwKF
k0jkn9TrVgSU1X16fNeYl/f85Lcul8wTVEyVattkqKJi2RIWkdaZQ830XyjwA3sqEf8AFXguAU9aSAbhMUpSj64WVpCiBDWk3zRHo1U5q6YGl83ZqAxvcsETO7hUzZa0
jK8WI0Jfp4y/UHR76TqWtJdYVBIA86uALWHFBXPDvw62DM8PyXpUDsCmHtD3SKfj0ArSjWw56Q6M4tc1/NlX0DKlvnM8n+ptRDr8hjYjEz51LuuEjiRPm5yAMD3Y9Fim
99ZU9Id4KkYj+jnRS1WcqYw04Jdn1U+lmod7j65idIgypb5zPJ/qbUQ6/IY2IxM+RTed1aINmcvXc1dxn53iEffWVPSHeCpGI/o50UtVnKkdMDlOOjbSWDK9L+0+ZXOW
MqW+czyf6m1EOvyGNiMTPp82z8mc4xvo/ifIQ1SuxU4zlCveq0vMQePGY8kWctn/jtKvCIlQomGtJPQ7U69T120E9qW/sl3BlyGZ2UDdiQ0q3spiFYvy+Pv09MoSIM3a
uKZtlku8RJr7deWQOcLJ/5CUKLDZITbOHVC/fNJRs3/cR8DEHiJMYqg0L/r7osPR926vh3JG4xuoqInGeszC1gbdgHGdO4Wip2Gvz4DtT5fn2/BX7sfDDnlThHnm6f6/
kefnPGs8VR+wQIXzQk4K39tQAID/ZEBTmOCatn0NPpkxikWQ0JFi0u9kRTfjtBLbbQT2pb+yXcGXIZnZQN2JDZmydC3BSCLVo7IMTE3swTT6ZOWUVHoWGUdC777Q8mvb
j+g69/0HrnvS5drhxr3rKm33DQj/lNbSEE6wiI4czO3zy188ZvtwkT8oOtm4DXGgCpGCtA8fMos25MTtkSOActXhYokrktB5KuxHlbHfduhPrgcUFhhXqG7dsvTg7zlJ
SV49H2EFcyRXWeFZ/lZr4k0wwmXrgGUkJ2MtbbQcispyuq5hUvj7LpsMst7nAArIgKY3HOKtNh3t9dyzixdUhFSERuGP2rX2IvF+hPhbUqIip4tmTuvt65r3ZpdTkk7G
wwFRIuLdJzqxHtOLo3sRZykiLl5ZI9/2QhjUZDs9y6787X7mRDDSBdwHSZpBxuL1l7Z3iYg4d7ED7hdBxRyz9+fb8Ffux8MOeVOEeebp/r8UlJqaSQrtllhli9K51Gin
j3ii/dj8aRWPmYpM2IRdnxNj0wEAQJhE5yXvpCIar9N6K8BRjUSxUCQf/0L/vZeM/nFraPTfQnFl5Uv9en5n3vPLXzxm+3CRPyg62bgNcaC3G496LNkNZXVUyhFi/Bno
t8Fu+K3JufLkWVUZjYCmCiVnRoZiJiPzO7VgPKg/H8svmx1RDesuhixDlBmeCcZHqwj+rT4/DmaLG1xKECpYXBq0sz601tSPxXNaFlXDmpR07ydzILVJPQetjWPt6rYT
CxbXqa3ZWJ2MYumZ1uB/KMF9ZHTMr2BGUMQZtw4mi02u9ysH4sn1wSjRHKQjQcUfHjOgfrDjF78VdZrzud53lPvEkTIqL2cYuFyCkQkoj4joLwt0dhi6dbks4+4legN0
tgS7lVXpG9F8pfSLbLf2u5PcMw8zH+qdvf5+bXa9Gib3bq+HckbjG6ioicZ6zMLWh18/rZe+XKMTl+Ck8SldB7iqaRIDuuEKVcdSm224n+mQieSRPmDxdNsR9S2zblAq
Tjfwxi04SDfYgv6MInXb9WyYAMoeIB9kDA5VRQX6CtN68bx4rHZkdPKhn8C2PZ3mkP2Bg6tjhRPDmKTS1tSsnNE8c6SdBQrQr5nvAy5j/1MO/hXWndELjKGGh0D1Rwu+
GLBdCnP8pwBkCWtywAVv0fTafQFLUmHtLSdJqaHXl7g3rnTx/bHq5YYMHPK/mY87sTkkWs6xmCoqgIPtWjt2LgxTWMgzrVOUD1RG5QSvmt8ROPh7wTmVNo4vejgt8cm1
qcEK5aAD4zfl68uEuuA1te6IhaLBv5nuzGmqbemaKL1t8fDRd4+3D8j/TuNxLmesuKq0GQ3MFrow3LsEfhVKFbKIleEFxHG30LysFECiMYNSkbmi8zwAwjTQDX+bW4DU
nBHo4GXk7hTrfeToAJZZv6BqGBboox/HuP5s7DxT45Hf1mf9TtdQhxTOjtaFTXoCy8w2K3btT5A6z6GEDCupP/a4ziBXSKCpe4VyfQrDEERLMB9dzMd/3j82eeZb0wF/
YCEDO62RezxMUXwpaZ/CUAXHU+VwCwruIe5duaNMTpGb3rhkJujd+zxRKpaRQHdYJhD/yW0mxoTtaMpCfHVkDAdOnkxrk5iqKoO/eSnO3CZSvXcUjedrFkjxhSxAcM28
fAGxopsBcL7c4aIPml8uGpAozbCng/jcNg4BEcjcYvLHN5d8rZaUuqFuigKX4NeXn/Wo2D4idFTnnM00HwuIL0tthOIIO3yJR+oDaBaCdDI8PtIDHHoA+MPE6d2rZh9I
PlKfNX4nnZoxIJDdlZpASvsry0g3lc3Qn+YigYl4cDwRfNzsiY1/y6S0io5+3uQ3138JmrxVKRKGUH2AsswEujBR1WA45RhRoSP34mlIIxBgQNTcfzPsZZw0CwnaJDyS
pOD+vhfPotimRnot4J/xmjujrlKhY5r/R7T2LVWxBxirVcg6zF0r2Ha1ICz2ZH3W2/bKtlshAIdjfLyduhFtRmFvKp26jUasCpzSJkHa3BXD4Ct2Eh3ncqKllvEOYcWK
FGiER4uStY9JGw3CGxUJFs7yYm6Q6qDTYyXB4pnjQiDPxt6JJqFQpS/EC1bt3kYgo09pxzG43rLtAHpLkcWsUBhCHQK4xURDw3EUU12B+rwXuKP4ozsLe+/g1d6aCPjZ
rr3/LxiT6C/jY/X0EdGh0UAQ5jbiwiRixlMvzCK8kkR2SmuDEvcF5K79O0l0fvnjxuBggLuaVKnbSa4XDz9NhWUvXig1hiXyhDj94sIVZvggNJBM7yEuRr3l4qQaiC6P
YL3vMpjZA/eO2aDmjv68BcY901kc+cg0lBAWS3a1nIxhcI52G2O0UtTUs+pifymxk20HBUCYrFIEDuU7IJdCC+6IhaLBv5nuzGmqbemaKL2mr/3Ygz98uhc2XOMazwV0
e+fbAXaxZ9iWHpsYcbumnrPpghZrWT8PUVSIsoCFDB4TOMkfevkT+jsq9nBfkGI3UM8UI7BbcyN1G1xCFI3kbM/G3okmoVClL8QLVu3eRiAMjE3FtRv4C98+Gxfp0bpy
TmqpmvEM2Eaf4ND0t4WctwfJUWQaHgbFmYkzumy43DJLxHEfQ7gaLecsIsZvKe9D6rfnoswjN8PSh6SrzG2Jse3I3DKhEz7Atndj2Yj9C+ZD1lY5XTCFIyT7Hfe5t6sf
+bWo0UQvT2k0KtnyjGO9e6wwrrUK+CD3SUnLyMJVAUORcZvO+f/mfiWEUUIcBRI4XYFDeGDP4lSqzbcngYePCrBKhq+RcDc4dlUb+zh5sJtpI6r4PyN9BeNoO7vrJLSD
qjSl1c9v4U9LlA9DSeSxx9mj1Z8PwNu7uGFYLRvffDq5PrzO5MHhv7yh4kU+3OOhNrJ6lrsg0Ck2mrxdU49Dmaz7uVXIdogDAfpLJFSILE1ibuDieN6/6YLGJ2h3d8yS
EhuZjB36cnGzTSWjV13/ReSSeaufaPR0920teFOCb/CwJ3PNQ5IEFdb1VPdlSzbqrPIz9vP821YId2dnvu/911K3BJgpWT/bhvqrFVsWdpvReobea4V5WWwi8rl/Jxix
wNnwaEFBwY3J1JwACLMKJFzzsg5NyAtJpOhm36VgeNT2aIiH2vU54dNzlZjclQCFdHhWalG201yHmCBg6aUXdg9yCdOp0JZ2ErFTzVrw9mG8KrU5au8kYFEBP5GN92N1
AsX5xNAIj8hqSJ9/7e0H2I8QT71txe53CDsAdux9N3DRX9xNckOho/wcuw4mO+qs1Da5itDcdyYKWb7xLn4sRtmj1Z8PwNu7uGFYLRvffDq5PrzO5MHhv7yh4kU+3OOh
ZAmdBP0SZikTQ84UGg8zbK0zZmRg+yKRqg5nCturMw462t5xgxqiQcRgul7a1+UQ926vh3JG4xuoqInGeszC1vbg0Mr/7ANJbipqnpv2VUQu908ParTNMcF6+W19fUuC
SENYJJyS87/ED3QCCgol9vZFRtnNtleiipT0f+M/Gwnc06WDAV/9SxBrpJuoMW0qnDweIHQgBAc2VKH2TBFKNVTJ9Nt3sYePVNxMb6oVaGAL5bzu3LDg7dwL6wMh7kQD
DQPTNgK9VmI6twbSTCtqgHMnM7yNJkFAQrVid3gEq4h4fNsJWMvdUtypo2GsgUU9LqivA8C4e0jbHa/6F2OFjgWX1I9dam64J3eVrgsJt6XI5lam4UvfsoAoOMUpGUiU
k5q1YXZWKOWU4DMtVTt5knK6rmFS+Psumwyy3ucACsgGdgwia9kHjjmNOPcQDz4Cyit2cSBiamduUlN4azkFNftjHrygFJhbTc25zuXOPGei6aqHqoAlNyCGcLLRdSSm
1IHMg1bw8M47SJKpBpC1qdtHTAz99j6xVxQCsR9QIOhwo8LTIDqERRXmp8D7YFV++J9h+KovGBMCYQa/Mj5O92wTSUmZfLWhMh4pvXC6eqVMghJU3ejFkTq7t/Tao4lQ
OQn+z27saTsf5/vBGJysxuzq3i0v5oTBznKpd2ZNL9FdRokC9Xhw5jNpwDHa3JWeLmKRiI2lIu7X97POMWrj63B7O6nB2ox94EkPd/bndkljHVakkbtYP8iLpG2slYx4
IjE1GaB+QnvN5t/w7sK8yrAOE9d7RIlxF2gY14AyCN93w2TA4y42PqbcFGgkjWQoF3N2vIhQOOY+cHZuVJ7r9ezq3i0v5oTBznKpd2ZNL9GApjcc4q02He313LOLF1SE
WAX0aSq8jdPnfYofg3WoHeYz7hBGDnzUNDDnpx9Sk10Pwu3/KS3b5q1rsUYSHUBtBvJdWrSxDRR+mW3y/C1/c7/ndwKYjnFyMreRiLYsnBVME16yqj1uK5GKgQI5L2ig
6OTVdnE2FyDiiztZEhE9upvYE2HnlNCT5vyDAgXs0Wmlgd/ns1d6GvIejMzwtSOemA/1nVNH0BKbY/LPFewctFBPVeKeDxANZj2j6qnbEQYcWdHPYxB18uMkj1Emgh2F
pDAixgPdhmk/Wm6tR3wtrCJAT/u5OTFKiKxQOL8MbZQXc3a8iFA45j5wdm5Unuv17OreLS/mhMHOcql3Zk0v0Q7f6diZ6LcPrbzrI1dj4T2+JG6zzXZift5o3lAtSV8x
kJe0dRu9ydSsdAOeehmyjliUPD+CIMfmbo36wMxz9OoNoLFGfnLasQcS/2kzJmqLU89LEFx9zFW7Vd3Gc9B5SogWwAkK+/H9qs1RP6cAm0NvZz8WHCAWbvpxrKsuEkA/
HsNKajPJSRSSeLFLCuPZoehA1A7NfA8K4wOiKxijzEAujnbpEEqNMe89IsafrMdU3lEV+b8hPgpSuzHm1Xor608iUDKGm8k2hmfx3N+Mve/EmBPSk0KCZ5KTVBLjAZeB
2OQFJmi+WpHEvJJYCXSZC8c40kxf+lZn34bO1gpWUTs4HvYqPtsFWUsGY+tOxjq2Bh1PIIfiZHW+/KBS0qKlmTYHXYgL+ycDuhVAjc2Hz24j+Oiii3Ru+r5VVAzj0K4g
kZv9eNh/USRGefgU7ZZkWnfmBlNbbXFEUU0A3QjxZGypke42a8avDa8r8kKYOYu98JqPLoDmHTjf2KTdqdArus3OqvbosFkAM/spQ1QrRbK3cJewEEjC4xGqg15w2DYa
dJuBBBvZlSde3VhOTgDmf5ZMNnTDV+oNJU03qZ+q+m0LAcaxFaqpJcQFqlQThIyLlSXZ8lPw63vBEw3Zv4b/m7s6U0YwUafWbFP5VK8D8Ywk8Ks9+UX76NA03Bw7NDhC
IjE1GaB+QnvN5t/w7sK8ykgeo58QewtOkdJuLkdnIrK1wnUPgJAzp14pKRNdNFIzLo526RBKjTHvPSLGn6zHVHTkBpTX52Q/OHkwyWCxAIpba59b/oVzuDVYnVbbO+Na
8kzNwQjwzW2EAnb/ZlcBCBYOlIKWRk0iwdce+u7eASVi2RIWkdaZQ830XyjwA3sq2en6PawlOeQRl6jfm6HlEDZdRNnLhs1TrUXxQv6suIFIHqOfEHsLTpHSbi5HZyKy
n2JTt1K8o1GaQxJcLS1s6CkINysCNi2aVp7J9/SQ+vx05AaU1+dkPzh5MMlgsQCKI/jooot0bvq+VVQM49CuIHCpWuR9dvAnnbD44tpGmdejI6li53XdjbsgT2kH9zVE
6yn4Ac0ibG7qLYWTTOs7hmPimyZJR/F9W9o3plNNX5HkZTcJx+Hiux7bPzSud6po8aueeDpm6fRHb1mn2YrYv4ZOjDhxYt7DFVkUIClERxWLJ2V2PvCiEGEO+KqrUptQ
UsamBW664by2UR9xsC/wDk+mf2XkDDhoLnYUixGk1goYACG4zY2L2h/IN9NrIY8u/qwfej6WAbjCFduvUmrBzjs+FcowHIPWZY/nMBcBQ17aBI00E4vqV3iBhu1KHnZb
pqfXqSphjQUZpSZjH4ygfdILvtLImYKbqdQNjKCXwWXwyZMGKvL9+243Bu1zLuCVSgU4J6QVl4dgW9yvUOfSrvmJBPFab9sxTnVJR1xte+uFfoGVKfBs5ERgx8BJxRct
rqOeo4ZWDeA39MOVfY5CJwA8zi0SMruJiw3m4wuAjfwVMSVqBo4PMDvpgfn4VS0nyOZWpuFL37KAKDjFKRlIlFgF9GkqvI3T532KH4N1qB0SJHaANvR3/LgKNPs9OH+K
oUk7QN5ig+UOJlL1iiuyrXwU+hYpRceB7z/UJJOvGyU24qMHjgPU2YrwJvRG1q0iUIONXohdQEDDO41sKex/CXGJ/PSrLUD/aS8BPWt6qlHHtHmcuuE1/VWVkZoMFzuA
92+dDBjc/sidIYyhPc5dbDcR2bGaAphglWdtQgQd+BiNU8AYlQLbJRoC+ELOKz65KsAfj7e2JmxOKlB2cFMV9usqO854CHc5b+zO9zSvCUdvhr0TysuYj1ESI56q74VR
u7REVWz1WCUOyfLLtPq78MNmc3UFc0W3JT0qrdPVXpqCBIaHYy++VRbmWaj9V/C0YDIoOskvpD8f2VdX7ATzAXn0igDDW37Kj2mTOd+C979h1X0MUNJAUMXpzihsz64Q
pXCxEq6m/vLjnUZdXviGar2HGGrg6lVU42mlYd9Dyw7bmNjAg1IYfBpCGrbKiFQk5JaCFA8+rKzT1wDrgyuZILGrzXUeizbA6eo+Jdve5G0GJwAmnLt895XVsDUje9pT
dOQGlNfnZD84eTDJYLEAikLfbDIkI18td6LDxdz6PITpZV+1WmjQoGBzfwGyUgwjevG8eKx2ZHTyoZ/Atj2d5ilmU6FgFCsxKFO6qu89E+euFlaQogQ1pN80R6NVOaum
H7unhdz2ETatGCF1FZpdqWLZEhaR1plDzfRfKPADeypOY37RgNcCNqybcazwwQeP7xNsfSnawPp0418jdqIPWDbIb3iGmbxVtCwjSG7x5kmYD/WdU0fQEptj8s8V7By0
itZyVmPh49FOMZXHVxTJFiEtpyJzxUvTubbO+dNMWvqJinw7RaFES2kiTfY1oQuesavNdR6LNsDp6j4l297kbYeRSVl6pziYeeOgHr72WiohLacic8VL07m2zvnTTFr6
ZjWTqzv6NHt5VmFVVLUfPrGrzXUeizbA6eo+Jdve5G1bOMEsfMjm8cjUM7D6CFHTIS2nInPFS9O5ts7500xa+tGmmF5/EFnTeb3/+cSPB0CkMCLGA92GaT9abq1HfC2s
PPA25TUymcMBpmZ1eEtPmlUiSHheRHfaUEecBpmAfRsh4iDxhl2dMDF4/Joeu7/NgcN7JPqxTnvFSUXRAumfgGRJJY4rk7InR/dwo4V7KRDkkR2fh7tsFEruRd7sriOG
ZizVc2/sA3Fp2ONaG7TyaaxnyweAEIWB5pEjjXg/Fxu6MqrstvmLGHlwb4q2xjYLBEYvZHt5fFBIYrFmathuaWuX659e9S8wh3pIrLXQHY2Jinw7RaFES2kiTfY1oQue
/ef8LckCM5LbZZLZX6BZ9cKj8OQiS2FFlkSpJs14bu9rl+ufXvUvMId6SKy10B2N0aaYXn8QWdN5vf/5xI8HQLnpQCE3du/nk1/NKa4qnhpGQ+qaVcCXydXFR7rYwhH/
nBC0CtQ5RXrX4R2gqp7v8+Y98ET2cvOxUdpkx9P8ixib2BNh55TQk+b8gwIF7NFpDdJaeiYYT+/soK7C8H5Reb+5nwkNVAvK63x1Hvsgeg2iB+ev5jfjn/w9ly/Qtlz0
c9WkkJWIV01hY4Y8C3EhzvifYfiqLxgTAmEGvzI+Tvc9E1ca94Zn1chmhAX8xG/mms6HN3nXMcCrWnmM2pYlZA+/OYdSDnfU+kHX609y58CKd/kWmsO/mBRbVZuXwvIh
dJuBBBvZlSde3VhOTgDmf/9oL/xtezT932VL+4B8sj/zFbpJ9hugDLjhBGW8XbIDwBzToZTWGP1y/HEvRxdUijh/LReaSZfenu3EPqRWe1Vz85KGOCdgMGccuMhJHaqR
J0eFsrECAtNGgYsA3kWFmUzaqnomSE243HgRBC6f/8MPvzmHUg531PpB1+tPcufAXNeGZgOExapMp94j6zw2hhCJLOS+HkbD+vejgUAUYcHmM+4QRg581DQw56cfUpNd
3A5qwQFFIaW2Y7QQU3B3nYDyZpbUbr8X0o/Xxa8ChHSFgvjVN0Fwaf5Uj0i2kl7b3vc9aqxMGeFpaENZyuJ9gMiBh+sSVkSotw9/mLNYJRESu025vVa9hZocinh9GTqF
LmKRiI2lIu7X97POMWrj6+A3RLn8lVGE4F4C9nz6SohPpn9l5Aw4aC52FIsRpNYKGAAhuM2Ni9ofyDfTayGPLk1p2SBAiUvHVJs7cO4xDkww7xWzt/i+oKWQ2eSI750v
BPsTV2DO5G1+A76aHw9pt8rvtEHogS2pU5DYQ0Eey3Fv8a9hcwu4qBfQ/TlOtZ45p9ykIgsELZId1ziqgCtFLy5ikYiNpSLu1/ezzjFq4+u34k8tJOqm39cy11aZ1jF0
7e8sZ1546VA9xUq29zitjgvl4CRvee3fbfkiEGEky8Io4BMBS1zRlrmw0MbCS1qM11vSeeC7XaXAzNbI5NUvhTA32+5ElRpQ8Yb9eKAEp6Hgpv1wB2tTEYClLqkw6I83
gR89AYsTf8d0A+k0IZ1fvo6S6doZhnSru7HiPnfAhzz4bPUdwbfNJmfscTn1LwuA/K76Y/e3hztaNVwcJaZD/NaajgYlQmKJf7Vn1YLUc/IHTp5Ma5OYqiqDv3kpztwm
JicR1B+th3WGmEbbRVcd7LU1XCK1P69770bfwFjPgey78e3TAh9CJZAUn0SjTnR1L5iuiJZcD8qjBtX/DDVUf0g3ZTPo/GDb6GC2Tm7XjWw7mS2siSkg3PsKZ87iqaDV
AeRVHpAfyRIEq1+RAVJxBRgokqHZFqEG2jeSf2KZOHDVPvjBXLwqbga8rKAlAGQXyZgKsi0LVf0exPgNljCxfdiTHw1QYIZsEsjtb5s/HECq1Mvat+wBVPBigc7GGi2p
QBI0WPWajEWouw+lVttrCf0SgoWN8AzQkku/gpsrcRCuVMQBA4ckrMQJuQ+5MQevQAgsmC3yMhapbscu7FUOzC/Ye2m+1K1rTCM/Sx1cFmUi6LU4O2yBGY6+nCBQ951s
HS5cmKN6TL+iqZDlUBww4sN1pg+7u/FxKycvfaI4BafRVj3JhMLoX/hkOShYRAa64jpQXBePODbs+fWVKLbdkiGFgCpA/Rl1Op/wCj8vJzGO649+od01MrV7I4rCvR5D
LDq6p/zwnp9QjYrKzg4GoRor6viYTSWeHGiQ0j7yDsGtNnSHw0I/6Z8YpUuXfLnEEKLv67Eyv7E3xyBPJRpPQK5Zc5ESs/QgDOV79WJieJrAJLN88NtXm5A8De8SirGP
yilbRjgrQzENrHAhaymo4JNvIxsKFxgDrTMvK46g/H6Ictewa4ZeKSdk1JIPkg77DEh5QKFU/CXIgz+CmmqNu1MGbdr998LatKRdqaWqUU+20MsPQEyeet6lD90+kQQL
734+3XLH9xrdmXyIHVPJ43J1RGgwXUDIT8y34+BIdP88VBKqY1N6ftakiz58aviCGCiSodkWoQbaN5J/Ypk4cKW9yq+fuiB9rhKxy2IdsDS+wdjRb6cEIqQQWS5BsnCT
2JMfDVBghmwSyO1vmz8cQKarqEMUPlHcMB2ReEUo4qNYmiDgl9y+/utgMa1GZ+bgRus6giZdeL4Nzi/nM2eEKCq/lusFl0Q2OVjFpQOEBHZfZ7gT01MBBYJTl2bopP56
2fl+BZboq6Jj+yuQuCBQT7ZWRuHRbLjQtZev6tqOFCusq61IW8dB8QH4gDAr2zKbVJpranePBKnGut57Vohmv9bZY5eRoQPufQu6yvAQQ5EsHcJ8qau2y+yquv1pe+R3
H2HHR4G+1uGt1k6lGP8eibOorO18Tm0KicQQ+2js3qPcSaaPCEQPAg2us/tdH8+CCZad66hKdKVv2G+WbKV5eAECzNKnKgRh94tRLy0YPfbz2T7/XnbKPisAgfcaj2v9
3dOhQmTGVjVJy+34k1dDFNGYIFk9UIRxQmlOnyu7smUOvZzH+BDX0LfWG8qhn5wJhx+va5f+Ha/AQKd7XWalI3ULh9UY0VJ3jewIKPpNoniH3dtAyVMB86Qtj44RYTR5
xw/wjDeDz2yjIOY/ugfYVyXGyrNCEV9vXxQPhgzsFhu370m7+YNeGLEwtZxvgq6UaxsOi4gzOfR9dTXoDtVKAbci5HrqaGCDZ5ot72VHJ3VSZzKOzgXknFjxXTajY4va
AR1hf02R28FIue4rJxEjjuX6SRywSNkVhwlYAUMhVFyIctewa4ZeKSdk1JIPkg77BErmrofzi10WUeKbZmHUyRiledl4MdTl7KsoaUs25ny20MsPQEyeet6lD90+kQQL
CeQbnzCF7HxRs+yAbiK/JN3kDi55dxwco2pxeyQ8vxxlJmDij5o1QrpYZexj9ANY2fPmCOELYyU099nkxnMaJ6XMlmELsz3g33UAVm/fOkc9ggpbxwouL+wZUPvWfFV4
HeSlW7YxqJZWHBAps8dYxTbPlWEY9LyY5vK3BOKIBQdPebI2ZySD9Nc7UcZbpk5A2Qg/dGZeCOxfn2W/BwK2qqnCIx3zDZRLt6iqJsj/P7F/QXQAldk/itQXYx4BVOdV
zbUf4VH0lzOqiTmsWodQdX5wu/Y1vkEbxK1A3sNb6n5uE0WJheCm7TzBeX1GAn40WBPhtAnhV9zG0NW6XQeBmx+mjcLQt9SHs7WRz5x+hd5D7DTU4kl8qHU3ktAHrrzY
GkRkiy9VfuvuefHkfgRAVr8ZYoZT8nonSHBTTRv9D+cRIhoeAzs+SCwHgirDqiJeZVrVQlBJ71+7GacwSNqOQFN4GkoikVmxVk7vu1qoDXAV3PjIjy8Lqf7W9Kk9xA8Z
LGkW1xIh+Sq25ktZhNzdDJDqmZafgw82axBDkXHlkZlL15pyfNFYvN3gaqQQjGX8WorFZiZ2n3xSQOOaTQ1IECOoV01L7+igawnbk4+zTYap6JZ5JhtAwfU+PTnVDnE3
3vc9aqxMGeFpaENZyuJ9gMGeO5rDRrozkiAtaZXkMxM9mU4MCmF5C8slrQDO8P862RSRGFSm7XHFhiZdlmAk7VGeIboSA7tdsu7HNPlpNojXyssDw0aVGHPwjj8DEved
ogfnr+Y345/8PZcv0LZc9NxV/e/f9+p5b1RiAkaNwLEybaDR38O6jBbNd90LZdbz2xDCzfjQZp4kwAcvN9bD9aieHbaKHgJOkYP4NUelWGtCDY6kpPPo85HB198p+T1V
8Q3qtGTqdbopCys720elHjGusBPWsGCGmU/Ys5G4QvekMCLGA92GaT9abq1HfC2sdQZGzlnqrvykaRT8x7SiJwg3LPgoRV/dXxuq4t6hNVfzxrVqIbLm8jGOYKeX8weA
/e9qPv5HYAN+nGJsjshrtbdWVX9ZfJrAi9ohaId6Skfdn61KE6lRri0QqaV6/H+8sRlFyHexUL8rAeqW5h0Hv5gt3APP0LRDodn0wACxTtoe8TAkIeHvsJg2vu/BwVsC
TBNesqo9biuRioECOS9ooOsp+AHNImxu6i2Fk0zrO4bbEMLN+NBmniTABy831sP1qJ4dtooeAk6Rg/g1R6VYa/OP4rxMx2SMOcNT24JnUJUg/M+RkNBRiovharMAYzTi
XO7hHnk/duC2aVOtdfWehhSIrVmL528za633k7aJ6WgtKa2m2zfMwXWoCkAXTqs9zc6q9uiwWQAz+ylDVCtFsjKNsoxM3ugd1ghXhRcFU51Q4UnBkDIrATBm7se0jqV8
eednrdt/LyamiZGxjLCYBZ3BdJnlU6ljxZYuyaLmBM2olGVKtK/6ceVvqkGCMmBVf3FosPuw9is4+zcXCkluQSHiIPGGXZ0wMXj8mh67v83rgVEHGQSn7Ip5lV8y037H
IjE1GaB+QnvN5t/w7sK8yu0uEXmWTy1Uj4Sehymt/kk+mxrRdmF7/SkuaV6ecLEayRMiSe4SSzLhZyDJ1nF062cx7u7pVLuFbj0TkJTNNh1Fjxk1tag1Wd31LRm8W/Zv
xJgT0pNCgmeSk1QS4wGXgdjkBSZovlqRxLySWAl0mQurp4qJIoTFDKJ36wgHFvXLiOaAGLHBYLQOWRd0k/mDFh0PO8KM1PvuLY2mOQA86bwVjoG92xmURnHy+7JLYLFX
qVu6MnaBCMysuW8+bF32tJCXtHUbvcnUrHQDnnoZso6psBCPpIiRstLkWacvgRhhZOfDb0YOZlyjO4u7mVZnNtuo2yo/+aX8tsJvmrERPgGxqOoZyMjylAKYSq/suwz8
t6HAN9xqW/uMNf48f3tlQAmMOkXoYpEqVjJ1Hm+f7+CDnxFpSso9Hvzsr5CT+GPrqJRlSrSv+nHlb6pBgjJgVUNhsPXtsBg9YLwHMMogcFqApjcc4q02He313LOLF1SE
EIks5L4eRsP696OBQBRhwYTWzJ1ix1z9Upge/PMAbFfIUp4yrsrkjJK4f9NGSXWbgwwG8EDk7Cl5AT+DxOWGqByg0qMYOVHvhcRkHespiWwJjDpF6GKRKlYydR5vn+/g
4q/B8O80x+zAmiatI8gfhjhdotvHM3Hl8PcGloeIc7W+Dqj6M/Y3HZQwCSGDBd5oRY8ZNbWoNVnd9S0ZvFv2b8SYE9KTQoJnkpNUEuMBl4E8nNYXyqVPZqEFf4XvIdWz
/qUOQozTq7BIjSo9+H7/jMAFbbMh+7gGgcPcRriXyTMyIy9TlPy2ztgdq+JE3IdX7xNsfSnawPp0418jdqIPWO5Ixz2QYxLoTNxG8a9iQJAdDzvCjNT77i2NpjkAPOm8
n+83wTskH1lykxhz1H/vvpZkwb/ybModsK1wu3TIjqLNzqr26LBZADP7KUNUK0WyUiceq8xVH02LYuL/+IDcoHSbgQQb2ZUnXt1YTk4A5n9BGTVRds6VVxR3GM5CiGha
MWxScFPMjG0YCA94qTzS0cHnWE4PreWfNzPnHtfYwK5S9W1RGEiwmdCf3wGm1egcqdg/ES9fgZ2zEBWqBUitgHuTbH+Vl+axKU5pa0FoxflMxDpIc6ReeYEafTpsO/9F
agUde7VkKYbduFXfBsRwId+qX1+C3d/yg0Ua/uxO/LnhJ/GtpzphEEFLy7/0nBZ9/ef8LckCM5LbZZLZX6BZ9VBPVeKeDxANZj2j6qnbEQbR37qdzHA/b9I3x6f/Xfm+
uelAITd27+eTX80priqeGiZ2t/dl1QE7c+41trwY7HwpZlOhYBQrMShTuqrvPRPniiQxJLYBSvfVhdxQV7Cs1LRPCkp/43Acxvo/6eHF7nG8h4ysVaR3QdQAUVYkSE8s
AJFUr0jPTolbfY9cNomqtPTBdhrXI7PA8rmjZvS6DBxVIkh4XkR32lBHnAaZgH0bSUP2zjGL8jG3FKXIb5VtJOmTqmSBnSVKUJ9LXE0hn2faQpz43inpORpmaQbkr86c
drgnvgXcBwgCyqD3o02iT+4+yRaGTjsQKfvtO/NqaXQpZlOhYBQrMShTuqrvPRPnowIgt2pPiqvh3jIrU4qVHd+D6AuiFsQKxLax/PWY0obS1EkGwlH2VzkDzinzp+fe
D5QEGnjXVrIkWcnLc6wZ1AzogvKA8YhbkJlvT2T4Iod05AaU1+dkPzh5MMlgsQCKx0EajygqHKu1LNxnvdFb5ullX7VaaNCgYHN/AbJSDCN2SmuDEvcF5K79O0l0fvnj
KWZToWAUKzEoU7qq7z0T54CmNxzirTYd7fXcs4sXVIRnWQPfesnhDC1kb3y1s0ITgKY3HOKtNh3t9dyzixdUhB+6rJ7Pt3a6Gzq/szqkCFtLbYTiCDt8iUfqA2gWgnQy
a/58hQYl3ACOQcN6kTFx/rHa+o9IVPcrQ1AjBb237HxGCl3aup4REy2st2qXhGSLIS2nInPFS9O5ts7500xa+jrVzWI1oz0pt9FVebxAzPWxGUXId7FQvysB6pbmHQe/
emqE6+X94cEoXB6TJqEjItlcncSww+aOX2bNs7ot896XtneJiDh3sQPuF0HFHLP36WVftVpo0KBgc38BslIMI/BnoLvndjdoEWY/rWC32AXZXJ3EsMPmjl9mzbO6LfPe
Ndg7Sl9U+HdABcSeZvHBxellX7VaaNCgYHN/AbJSDCM2/3KA2CWvy4qd7NHoP1Ds2VydxLDD5o5fZs2zui3z3gaMrZyQJZIQFGiR71ov40ZcJIfwPv+DTbn9rRre7BIh
3ZxRf6QF3YOhXQCMrdR0veSRHZ+Hu2wUSu5F3uyuI4ZmLNVzb+wDcWnY41obtPJpgoZB3ey9XjusyPBrT2fLsybjIKhhvpMgVz1f1e+NNnJ9GBwzb1kK3oKv+m2Z7UWF
a5frn171LzCHekistdAdjYPaegXL1y5CaQyzW19n2rjwyZMGKvL9+243Bu1zLuCVIg0Id7ITvclmF9+64ksOP95RFfm/IT4KUrsx5tV6K+uXtneJiDh3sQPuF0HFHLP3
be4K8eN451NU/m/gCn/VFf503FIPftV/+iFcCbjubPPeURX5vyE+ClK7MebVeivrBoytnJAlkhAUaJHvWi/jRtYAyM3X9pwa26LfldV+WcSpeCERDt5oi3A0ohoUGqLA
6ab9ur/IsxPHBJW83n3URkhHFgKj3Fec0eprTc0ferpVJyShl1AYf/0APj46DlsFYM19dYvShFdh13e+CmA7Of+IlgU8C/f9i2LWGgRenblrjkBAT4K9Fu0Qt/XM+emi
pg0Q1RIDKnn5somC71NhTG9nPxYcIBZu+nGsqy4SQD9a6uo2AVDUDZ+F4UCB6i7Gm9gTYeeU0JPm/IMCBezRabbYfOn9u/HnGp3rK1Z6NxlH6xOxSuYx0DATadgRE2i2
GKp73blVz3UUxxPs8JYt5gsyRqm7J/v4L4ai0AAOgS23i2idn+4+yAXWCD9twfyroAl+oNTCntrH5tLCT00/PsqIJtEmvYeBjKtfeWMCbYiYhx5OuEvGsFjraHC8F7Yd
gS+opxLiSXpl2kCJTQqWVhjH17LsBIppspxDOEufYY6PnUPjESU2NhaOO/IYMasgL2af1DWAun7Gw85NeirwLNOrBmC72/XO28Abm09BL+uoW+MxqHOlS1wWZAueZULm
1JHoxH329EaXlioiygG7DNvlNqXOaLJaYT5jp4ywZqAN83S09NvW3ZXdhkpqRvC6zFw/IBVbHmqBEctI/WPLcVRZCNpqQDF5E98Txa3mohVXzkrPveNS76UJhitwZ1mE
ynABcufwcDvjK4jpFBqKuH/7zyyXNeVKFOYZas+tsUiRW13IdN8VN9YgvT8aSjQpjvO9Bn3EeCLRjTylCkLRoSNGM+mLQRXWLPzbuq/GoT6O11S9M3vSgcRh4c6CG7Uj
iQNdQ+wyHwn2eONmuDAVmRYngJB9+tWKB4u8vHQ+yN0NoLFGfnLasQcS/2kzJmqLzw3c6nGRL4vAmsvOvoF69VgF9GkqvI3T532KH4N1qB2E+KPMVLEjfg7IoqFg6aFd
et/RbmBR1PBL9Lif8Wa5v+8USFSHYk+j/gGpyjxbV/KrUq4kn451RO+zDp7fUK1v6dPho+a6LpnUoMNiKAOqXV+IzxsCYSNFVs3PTomiy7X8uRTCCBDTsbBc0TWwqyTG
nqmJS6XafthndMSXIXTkjnSbgQQb2ZUnXt1YTk4A5n+jndzu02gOd1O6t2wkViyOY6xm03vAe4b/2ODdu0ZlJWSNvujCRsLrRe9Ukc5bPJSM15cTBBdEVpYggQ5it/o1
QEh+FXOZiQ2NdXcww0KYjDs+FcowHIPWZY/nMBcBQ16N7KLjPLBthmp7fW/lYRfK0F6dfF/yK5YFIFUbjSb6kGCsvds6uNQn3VyBx4GNCIuN7KLjPLBthmp7fW/lYRfK
a085ZTQz2kYtzsFA03PnEa8TOE+3HOMqEQ9Rt6W9sY3Pk5jZcLbEzv2Cb7qKeZ9S3vc9aqxMGeFpaENZyuJ9gKOd3O7TaA53U7q3bCRWLI7LttSU2NkBez0SkRpkw01h
nA2l+/VY4Oo8EUKZOL0FtTDvFbO3+L6gpZDZ5IjvnS8xfEo3/ZxGbgp+BkqL9J3WpbAKn1YBZh93MLSpuglKk4MMBvBA5OwpeQE/g8TlhqgdDzvCjNT77i2NpjkAPOm8
MXxKN/2cRm4KfgZKi/Sd1nb+W8+abV8ZIo2hlFvHtDzgczyaN0pMserNrJ0kpGToYKy92zq41CfdXIHHgY0Ii43souM8sG2Gant9b+VhF8oJ984gHBpEG4bY3DE7U0uH
QC5iUF2TCppOy3LYBNhGh9kUkRhUpu1xxYYmXZZgJO2ny/1EiXZ33MPiHQusEBog51MxdG89BlJDZ0EhK6Dge5h70bdx8ABstrIDx+wN0pEuYpGIjaUi7tf3s84xauPr
MXxKN/2cRm4KfgZKi/Sd1viq9yrdeb8D2PM+arBWkxSpW7oydoEIzKy5bz5sXfa0BfHKrlqMjn2lCcHNCbhNGAB6JDC5DeigV+GDYX1NMqhc73trIAXqsy9AlBm1CLuw
dJuBBBvZlSde3VhOTgDmf6Od3O7TaA53U7q3bCRWLI62rZTOmToWV6A+6/JyVpdLQ6jMrUk7F+b2ZjtvgP+iHmSNvujCRsLrRe9Ukc5bPJSM15cTBBdEVpYggQ5it/o1
ZnY/DGhhERg9Q+mgSdpcDnM+Rj3ITx+IhFxW0jrQWj4uYpGIjaUi7tf3s84xauPrMXxKN/2cRm4KfgZKi/Sd1grapZIMasuf0OdTuSHXRhbet0d1S3V8ak/PTedOmkfh
BfHKrlqMjn2lCcHNCbhNGEZ5sCGmQlItkl9LzLCNrKapBeJEaJwX3I3ujQmF3lhAyenEvXMtRiOCkuR1OvGXcIGKXU6Kwui6XPYvhz0oQS8PZto8pFkfR16UOuF+PFzW
0hwdUztih3Xp5igI3Ztl5C5t+XCQVidZkY6XmAAQ7P5ALmJQXZMKmk7LctgE2EaHfphmSvaqgov8aJB+sQ3X/afL/USJdnfcw+IdC6wQGiAJjrVRIGOS9lwkSV4/jQp0
HQ87wozU++4tjaY5ADzpvBGMeqKnkcTdJPlC4K3cF/E/4y+lnuANuGQYNi0mxR+hLmKRiI2lIu7X97POMWrj60Sd/pPAeo+qPunqc32L0SEHUvmfTHuM9rZy8H9dMrze
haY1QlSw67NwJWVP4ff0nRhXEIOgaNFowV+y24vbP7RQ4UnBkDIrATBm7se0jqV8AeCNkBwHeciB3o8z2E5HB07aJtzNZoqsyWn78KusZ9uDDAbwQOTsKXkBP4PE5Yao
MO8Vs7f4vqClkNnkiO+dLz1yMNER9E/mR1+nB3pPk5o8qX2myRqS3U4OYQG19Z7AyenEvXMtRiOCkuR1OvGXcJ3w17tq2TAEGbNGoN1iTbr6+/r/ObdigxX/6Zj4XLPD
INCra0ICeLYWqYC8KRGd3o9L14f/9NC7LgQWGL34V9sQiSzkvh5Gw/r3o4FAFGHBhPijzFSxI34OyKKhYOmhXeP+5vScjrvrjY/AxbSYX+TbwIiRBfqWlGJFwd9UmbNO
YM19dYvShFdh13e+CmA7OWJPsIEdyZr6j/5Ry198fJxaveUA/Eecg4c1faBp2Uxva45AQE+CvRbtELf1zPnpoojEvpq9hW7Ps8jdgVehnmpVqpHG6qDWHHBgkB7M0PcO
LmKRiI2lIu7X97POMWrj69sij8FNz0QBhB9NpqFCWqmpW7oydoEIzKy5bz5sXfa0/LkUwggQ07GwXNE1sKskxpa/mVl3WXewVWeWFQrWAAVPpn9l5Aw4aC52FIsRpNYK
MtkqkbzzQ+PdBonCeMYcderfSpepYV7pkiMqxiIm7gVShpIHg/AIpZ7VhUJ7hkw3BOu/Rvltd/hdf07jmjVfiqL+8sBAYnDeYAF5dFVjshI5s8kSv8aaJpf3MxyxvhmJ
jNrpVyXsPHTagFxhxNickVdiR8eWjBJwqz0zn2CpkadeHdBn+AA8OykQom5cW1eJZI2+6MJGwutF71SRzls8lLkzrWgY0rBnbp5pcxxuEbEtKa2m2zfMwXWoCkAXTqs9
1qzD1dIFuBDvxd4bVJM1ID9lybfms8MAPAIVDulRqxRrjkBAT4K9Fu0Qt/XM+emiYUedFKyEgYNpHVxExBZRZJvYE2HnlNCT5vyDAgXs0WkR82VL5f6cO3Pdm/wcFrZr
m9gTYeeU0JPm/IMCBezRaXPXZh+ASe5mRtV1aYQjhOyb2BNh55TQk+b8gwIF7NFpMcDcrS/rGEq01gip2YmxVr1kVCqlYRYZC07/5l5IFE4rRQPV9SFNuPBfOqrVkV3m
P1gDmwJmD1qmgbe1YadBdYHxegJ4bw+XvYot2cIrSOTnMD6wV4BX8AJtb6+lpLPc2oJwJ+eDbXCywK7GYYIVucJvx42rp0xpN+ypq1N76SM4rJ9PfFjqBAr0dBJrWC8E
rZY+XdSkH4lY6omSSWNTV25Tsjthtj/gbwosjjj649yLkil0UJwP4VVNvOw1v37Zq7OtzGL+nEsQfaoHtpD9HfXIkaNgSvgGkT3NvAYFid/m8UYhoo/lwxp2GL+KAEde
zxNRoGu/TrN43Rj/TvHfWVGi8K+QXQ+b0ucrpT9/ntOxObTs1TASgSSRUdEZG4HpzAfvXGnYjp5E0NJU6HLxet2k6x5ep+9bLcpMneNDrm0wxVPGaoJKHA0tAgxWGa1X
nyMFzk7W9pYBidOQOLFnfz2u5hk0Qpg12dl3+TlBb3VWhdEbZF/Bca8HSaF5jaWc+F7slNDh666277999I+ZZsJAG736e2UZAVErPh4/JHK4Q3sbS7bZy19jxiOpmQSi
ryyyTrEhwGy/OjZyLXFJfJojIO4XI4U6b0CalNo+B7OFc44CxSDF+l9etNZcUKBayogm0Sa9h4GMq195YwJtiIqvRXqa7Wc5R9gPXskyocPt6pn2/jqSV2eUIc/NYLqj
MMVTxmqCShwNLQIMVhmtVw9M0SnZF2rrkVweKfFl3ltU7jhnjDFOpUuW4x2zyGJm9L1Z4abt1n0J6bhciqrBdYbcjY6Fw88/jODx3NLiug9RovCvkF0Pm9LnK6U/f57T
hGm8aUChK8J7eVrLWBqbej2u5hk0Qpg12dl3+TlBb3Wl0ltMbU7fRAUmQXgkggXABBGg2U7Y8NtatL1SYWnXPUdlVDCQIyUXoYHE+YRIk6CJCuxhcJ/osFD5XNjIgNC+
AbKdSW73GHn1dB2EPYIcoEdsTxHSMe8UaREA9s/I8YEYAbNz5jpgCx9L6Kycwo00x9tGbtfJ0+NgePH15R+aY2ss21denOMorD5vT09/mJgaS1t24yH06NnxN5rCyLa6
osmpVpGfUL5CrAklLWXMb8c0v+qLr0tBGsbXFRRbBqHaVs9+q9EUfriZBvDEE48tGktbduMh9OjZ8Teawsi2uqLJqVaRn1C+QqwJJS1lzG/HNL/qi69LQRrG1xUUWwah
+g95P7urU9dWfniP+g400kqZxSgmLt/I2IGp1XcjXPoGmtf4hoTGN5lSJ5GhY51VrPwjnylPOCwYSBC8pMQjoZ3H8mDXduXrnqyEOSxv0u5j+4gqUBEw7adqR4d8Nhp7
rZY+XdSkH4lY6omSSWNTV/xtB/4H13mSABdNwiYFX/3wWtF3zxZmHwaQOJj6FhtsCXegWUHQf53gcMk0FUjRMSHDACtPy2seHoIKqFkVI7iySoPTebqlI8ZU9EuLj3/X
glWQ3ZOprivT4WSgcTW+9MJ4aVU78MKCa/37RhMQ4hNaPb+Oj5eEjNeQ7UZYBZxyuYoAMIH70MvNSkXkQ4itU3197f7reBoT7VlDw8Oo6BHe2DfolkiNM3wPtVD1H9Wy
Uwa2tuXz+7b82JjQFTsAcpAfwyN4pSx3pRzF/wf9mIPB3VLpC++ZQW+J4NOjqMzgmsmERYoybiOsutPrbhjvPUflkIOimGXaiNCPgc01B45HAtzFhnfzIxT6TKL57cyL
xT4STzbR2lbL1NDVomrnA97YN+iWSI0zfA+1UPUf1bJTBra25fP7tvzYmNAVOwByn4Vc53rHCwDs3LiptFptoOG8QD6WFf+7YdqwvOYj5qf8bQf+B9d5kgAXTcImBV/9
7T1gctS+ESQq+Irs9yEp2vLx9UMSOkxOZPgKPq14hXNRDdFxVUu6jx/wD8MnQU6xUwa2tuXz+7b82JjQFTsAconkO1wCQuan01rVdPMLnOJRnyr7LPfZJABZQQHMCp8G
vYjTV2Irypmn4h+e8n9pmAl3oFlB0H+d4HDJNBVI0TH/5/xcDMz/i7KO3GpHXRRo3tg36JZIjTN8D7VQ9R/VsrHzUxJonqzHVbWkK45+EorUZACCl+dU3B/TdLf9JLcf
aGJM4tcjmjsRh0FhjuWcbDd0apDA/S0VP07kUVxY2DJ3NhFJimsRasEAGHoikDVHveYdYbNDlTUX+I+7GG/qOn7V/6P8Xqbo5BqhLEPoPWxLa4nqT17ssjdZT3KAMJYO
q0cfpJH92WiRnbExuUhdwXVImY3Bns5qi0wTICFe5XcH9fFDOeMjTsIWgJI7zTJHAVJvjMBSzYP1kXfyxklFBOnm5i+2h/PiNvu3x3SUTuIl7YHFRa+1ICsx9FOFR1en
/iVXZfMJc2Vf6F4UPPiplG7eMe3EYjz5Hu0hu+LXbqhgxyzIFe49tSPH8PoqlosUkyjNbvtloOMTsWlhkUC+SmKtzd13zA19waE4qkTGPkKjMIgbMmsXNTEFKB1L2hBQ
44FI0w2yq6YYBW45G267+atiTXOZJ/hEE+0g/2OCcEiY+RIGDe/HkA8x0qstLUnvkI3WZHgsSzF30d1W+0gbAbeLaJ2f7j7IBdYIP23B/KtvJ8EHOsxmgaa9fXqGeKP+
YM1lbX8t9cOAIdFaTsmxUzbV513lc3/eEEYp5LP+NBEQI5EF21MS0A3jyhdqNlrKdas80Pl07g6X+LwdPfE1iVcMfg7MKEuG9uqYte+EzUMJkfW4eTfqdFPiz5blvX8Q
aj+m/cH9jYGxIw7xAleRhPjG1lzBACKiMrrnAGRyLA+9bxsJvRhj/ZWh/K+J464F6OZ+y/X4pfSa2yiUisez8sHTLsNA5k4/4Li662pz4hncD8/GBBhaBgkLK12fVWpR
97Os8B4Sz0X9SdyqUBwUcci0lAlQoH1vFmbNFm0hptPKiCbRJr2HgYyrX3ljAm2Iu7ZKCNBqHelcDrlU4jppFiGttWbL8KLF4TyeBF4m7briHj0rTxoZ6bRub8ATr+vm
YBgSdc14LnV1BqeUIPSNexVxtWrs+G8BZm4t3FdGZFM21edd5XN/3hBGKeSz/jQRECORBdtTEtAN48oXajZayrTUCosKEQhYZ66GoiCdZLqvhAD2fIjTUvUBvQ+21hgx
DX4RdxwrCZYXbQjet3UiV+uC1QeYDoMf8LJ0Le0kx04+EVjclhk5GMVNqGoHM7qC7X5JrRleX8h9cgBr3BfAUfGojDrhFZSMnBztdLb1ea9DG8FYtsToNw+ZZH2gkWrc
CZH1uHk36nRT4s+W5b1/EPnYtDGXlRlr/04bFvwXYYgn2XLG6/AEtCF3LozFA0YnakGXWJ03BTJcLJPi4sQoqD7oQTe0uF9GysgupuK51MtV0kdqSGBIaTKbOY5/IhLn
GEf5uu0A03kLix6vIdegDTwuQZJg5stv2Qpz+1M1aoojrC0+rz0wYE3o29HDFTT7LAG7skHSfdjoQLviPoAvcqQk4eicZw0l93JcA0Rpu/rEZo70YiobYs/LKyMeaiQF
VvgNP7CtWm13RpJCjd8RE3UxvVo1m/B4bkWg4ZdRSPqgGQSKaPwS2xNiuHKFL/W0pXn45MisM7uBU3jsjUj2INHq24dTdXF8K29xiRdqGFDqTNOM/+M/27+bPykHnA9a
GjR/Vb1/UBiGRQ6faR1kPVyAlh2gE5EaguARhpeEQtKKstG8wEoOo3xJkQF+czax8wYZ+mBN3x8ceCLXKpz+ROlD4vn2X29FxRhCyLMsB3ZGoSf5YVbFXzs8dbuv56I7
R+WQg6KYZdqI0I+BzTUHjkcC3MWGd/MjFPpMovntzIuxRjvAccxQNGa5OXawW062eQ35yujXoGyu4mG4OxdrQAHBMRZzoO+mucBBeWwcqCLrvK0lP3U6qWTYtOfJWQBq
uru6uQvXvmh4EkcizZa2N4KRXXh68gTmxo6mI3dtTi/eWEUz25MJw8INuAxv+cdwtKTwGhGAMnThi/rRMbVyvcW8nGuEK02yIiYQwuAhfp1y/brkB1mTVJP2dd/xaap8
9swyundbGyx67EbiXCt+/ehNoivL6TRqUOXQEhgoVpQJ5cwTgnGsuMdfziALZwEM7+2Gs/rUAQjk2+s0yaow+7wqtTlq7yRgUQE/kY33Y3UCxfnE0AiPyGpIn3/t7QfY
jxBPvW3F7ncIOwB27H03cHycT56N5Ze1c/eLQHSsUnDcpxjbTtEsgRBP5Z2W558CVBPdRzgd8Cqy36PCl4mpumiILTXY9HvSHGix38APSAyKLNE6ifXoxHRG7PTWCVhq
nD15WU/85ZHMBpTz9s9LoOvj6pRfZBUXNHvYUWd/y3JFdZaZKuOAvTCGbodrpqUIXsdZ6ecw0/sfGpi4BYupTEflkIOimGXaiNCPgc01B46DmHQ0ZXX1TugGODYmJHok
50QyuZfa95PP8tkbsPG2T7c/DJnozltBpMkWTghLfoSnghLxYk9jEMezhCSB4xmtXtz2fFacxULB5FejHsD+IdZ2PS8H36DETzePr5Q/YLkamnW3/x4T2hmCTlSFI3qc
j/+PTkimsSmbNd1yl61u1BA6ymrlcjnlPPtd8DroObzI82+pDXYNwTanO3Oj8gul/f9JfMJ7s5UwaxCAf9NlqqpmB/VKu7S+Ay0kh6oSkxvaVjQEbRJHgIp/VushHEr+
DioCI7UgVYHLr6fOo/PkpbcHymMc44U5n0IoH/V8Rolw4Dckfp0Mcp3KZNXnk3KRNb2rC8dNjwqOq3VQWYrrRbqzAlZCyjyA3gaiOymGBgoAcmBid61FsUikVpKpE1wa
MM06zAsD2tJ1Gn4dkASwNhceRvob4yKS9Z2rzE6YGpafjkzDkB17XP0lDom68b94UBshPJuMTd2M2ivSo15skcg20IZVbK+BlhmCvm2P2YvT4HESCMGcYwP6WEobOIz3
zKw91Zchd9ucxO5mTFxHHTdretrIXVC9obIhMTViULfB7dcVdqknwfMZWmvalfJO3LggGf4e5WVhC8+dvmFaeo4LzwAFl/1TNGWdpRt0dReIj6fOi3aEYDGwhDCdQvYC
zM9iOUhMpQfkqqt29+59jCOORHkO1AvBnrGY+mpUXr1sC/L/c3ht0sddO0N2y0MRO2gX8CZpmxZaS4vadhr50mI44bgmqUyjMWf5+5BwqrxiVfLkyAVo/t/GbVVwnt7y
GktbduMh9OjZ8Teawsi2urCfqgyOPw0jZI8tf28e07uaBW8JKAgVbGBbRtzWj9jXlp0ya//T30to7GiCAGfd1UPsNNTiSXyodTeS0AeuvNhTkP+JxSy35Knmph/GAmXD
nvyRvb2wRyOezwR2C1gekbPqBxDWpBRQwqHMOas8sEe3zerYH2RS2Jkm93yw39WLde74bP3BwMGef0SO2x9PYFl0FcKzx0/8nehGztSzdV/KhBAjxi3pdc2uUvSGAaly
04V5i6yPWCr6StxTQusX5K16QhvXQaSUThXAHLbZr/L3VDMt72DH+RwndyeHppHnsYba/A9KhtksiXnmWuYC1JpWIsGjs3o3bkTE70InA3ATPL9tJrRz0+bGR1nVlCxP
cVyNcHUnn2MDVEUKK5fJjn4chygdohyDQwHja4r4EkyTjIDJ9yyt7VR8MCH7E6ipuyKxVlnDOK1gOSDNLCv7+5hy9p1Vv7b8HCK4cxENliufyh4Rg2UAQarJreDFUlYY
s3PyN9Pzq0/lHyYTJptC7uQhUxa4/BtrD3hxEZm3mjQOyX5tkj3uhVdQr2tEOd0ACryFKeIizi1d+xLp2JCIZjL1AYMT6G+idwlbq6QyaChEx7K/Pw3eUGB4J/eu8i2T
aT6P5vnV/h4zESfyplVVqclf8dLogWPZSlaA9Fe+2cC3dIc9eMWKvDUU2CIpyqudNs+VYRj0vJjm8rcE4ogFB/xtB/4H13mSABdNwiYFX/0w/pirxKQJaLfU9BD97kgH
QyfhrU0PeRzyoz5dxnW//SL88fXX64XZ6fOK1BajVWqEXaPbPtx/iFOnpzFVOzaGXOOfMnnf5wj2BNKKXFKlUTqOYh0w6moENJ4VUEafB+SqIrud+SQ9WQvCNDXr90gs
bnWZCaCR38HAKDIhOHYCec1lm4RfkcmglbM2UNxREk5wuLjbWcUYGaXBVjo1VdHuIRMgbScZOxfiFB3kYaQbW91eEdQxAWBp8ltE8tpMGBZOP2//N1lipwsONOtvjE+p
WJYRH93pGv2h38K8bAoTwseC0xVwYzFqZcKNOgk0dfvVdCWvelf1nnAHZOUIH8mKosmpVpGfUL5CrAklLWXMb8c0v+qLr0tBGsbXFRRbBqElL6Q094C7QWuS2ftzODNC
MP6Yq8SkCWi31PQQ/e5IB0mvVB4cIBVQrixfEMjBKCXk+9YRHR3vgBK2ipDuixzF9jFihva3m/c0ndrYV8fZbnoLMUfw1961jdGoC6Tyyi1vmTYzJaSMYPpDI2DjeiBt
263jccclDxFTRVsWwULSlWUb0QTCXT3Yq+k7JeGpfp/wMxGCtH+47RTapLD5+rndGH2dHyr+W1urwYSQykNaGCbcSmfOnMZYy6u4h23MYsu72cR/c9hpMdwlqjwnIul3
sENFyX4Ec69JkDnI1PUL7nkN+cro16BsruJhuDsXa0A2E5zNats00BTgwaXvOWHjYe/SIvOjWfDX6gM4DvuoYesuAuF8ISZB3FLQoISiDo/A4M7FLI8JtKt3N0itsq6Q
Dw8rCY8PmFaDe4eDhdGFt7kULWc2S0UV7qGVLOwt7BrwLV43DvnEy8LKh0whZHkP5qcdwX4ydllxjnSN5dUTxiHfgBLxc6rJUuhIqvpnksnBsXKDv4H9ZAI5skrDJu2O
wZztWdD2W0/4ZBmfF4luQ3fa+UL7+2D3fQJ1x12t8O3YR6ZuFNOkT4s2JpRh04aai6mizFJaAxxjUBw9w/5oYpXkv6fxzC6uJCJofLxcNisV/4hIpgehjvBZNuL5hoRr
bgnceyGlN4M7It+lqQN0qTt6BKBMz8trhQtyHFsVm0GI1e11t81KkOrNkxSJZeeIfAGdjTBVy/9EIYvAm3miQsN50+svQH/rV6nVziPgsVlnQ7rrr0rQVNMWgJeli35g
RbSdtGmDJmDApG/7Tb0SYKu8Hl7RqDqGZRfb8Hm8u513KCYR0wg+icWdTfkNLcg0ihw86LSI4toObnc9v+z5J+Q3W5tPmYle1svffA6miuCsMCkKzDP5EIzivt9262Aw
R6l7Z3Pbv+zIzJOndgI5iUMlfMQrboub9l5+bNVKJM7kEOAqXDSyZNx1/U8iZNH/syAEmczvnnriieN0QL2VEKz8I58pTzgsGEgQvKTEI6E3t5+TuWAKfp/rdnIJQqNl
H2JvWVz43qYSJiHxFiFWOeCq1WU6agNdZrjdoubD4eYEvtgxrJTSlK+5JOQu0DTvp4HuQwEcRqSylMNwOyrIdMufWkoPtGwrCXnkvatqUumvi9Z2GnHrP1JT6ALG12V/
BH8FNa+VjFskXjnrh9FdrmU3tpva7Z4bmv00tLXZ+KT01RRVHzTIWO+VP4bUHWnCRRpprXk8uOeGTAgVJepFhoIRj66JR476hS69hiptybP2IVdqnM2Rwk6bc0xAW+Vm
mSaFflcRBvmjRCcTnXbPkVzlAjVr/PVmteKgTRzjE9RoYkzi1yOaOxGHQWGO5Zxs8FamG5kSfLunitpqwocVl+BTWNfV0Iqk9BFptLGHAJtstjCKkM+xCSBCLW+QJwJB
JSO9JxQIGrCSi0KdLaLVmvuO+wJaU5qXCxm6rRIPWLCpEjCl8Fwlg6WJzlW2u4D6+gmtLNk7JGwPq8rJc5scXuP0UW4sBNm0WDfm4WAPhmLI4B8man6auX0KIktB1n3e
vUC+KvZJQLLdzdijzt0hvbam0BilCcAE3WWjMO61Wi7gixwZnqxwd9LqKhTbDCzEaGJM4tcjmjsRh0FhjuWcbK4wZI9H63KJJYWfJKL25x4OSKhefUJ2vsuZv8uSbgpX
M2KkMpDRcO9OBV90VTNy8NIB9lFM2vLumGNIgvtIeFKjMIgbMmsXNTEFKB1L2hBQ7f09kXvdEMgXnIJ6QR/8DMtNMSB4CV1fcoIEsMntlNgjBRSSZJiK3ckzksm0zLiC
1qviWqzmc4NEq+X7rl5wUmHQ/qzG0PH8TzZL24IBLRGBil1OisLoulz2L4c9KEEvWhdxaNCiCa8Cgaynhi78X9Y5cp567Onf/0eHrLJb+F9q6cm8AtldmUObA7ZIXHWD
y00xIHgJXV9yggSwye2U2DIEQL3i7EmRYdgKUTJtnOyASAunzu1/jdhEo/d9tbiNGWu2zMGtnDVb1O2RFokdpIq4Mhw0YM+acgBjjwyTrc6E/nCHqt+GYqnjPSekfhq7
YR+sJ7FmthJuCVbE4ejPAXrgWvNl84U2r9GQSoD6to4ornLAvRjLYhxTqOcC6yqhf3UqMeyyhYJ8snpwf1njBnJDOauG79MSOydJE+fNSSuBil1OisLoulz2L4c9KEEv
HS5r8MdgxwQ48JpgvjcGEe4hpGfnrbJIBw3Pl+DxPssBG3Huf9CQj8SYa8/jVWR7sKjr2Js3azzwFpK7G09FYhS9WtAmO6K8vF3u7AXjgAoeYC+plEErOOErpRo7ZwAA
64LVB5gOgx/wsnQt7STHTnhZZoJXuMZgrh8KCiR7c6vt/Jvji24VGRrXgygsyAbTGLMWplerIeDgoSLkNng47mGk67ttKIFh2wAz4JtzVPyG0Z1gLWB7sNcaqPOT3kPM
Cp83PqArBDl3e8og+SdFS2d1d0687Ezp8WKkC8D30aHGPKc67M3ZHyJvFGKCE/25yZrQxiN31rdpEzA64G7E5pdLzWSp0Y4IwEK1WE98wK6WItGLTr15OZnMnJS27+Ox
3TOXUZrk1w/ewWWyy3EXlfZbsBIAfMXXZeGLEdTp79POrU4wARdCx3/KO8GTJn3edf9l/7ochgSH6rNsr7pdb9pltxHR6RvagJp62OMUMpVNGb3A6EM0466t4CTV3uha
UsnYNYhQnjiTnXPg78tlxXLXmQUJD4BIIiQFIRtXOagZwt2+am9dznvsqySdD9hC2xkwok7R47tklYdUY3e8cdP2SxjX44TVx3aCleo95bNoDKLvHg2DwgP1jOTJXO8s
7HSN5GWWVuO0hHtgOEbF0IDPtLFBe3d9rj0Tm9jaGDtRLszihsD4W7cRVrBAsSfJp7NzkcCSdEsfhqathU9BStf7XmDY1V9YtOx7X0/Mc9YW2DBbx/d89GhEqzYiApvX
n0CMPFunT42YCvZXlb84ZuC0DlhMpbbSffwEXBxiuFExlrhpKcSu0JohiCtH+qEHz+r4lwvOS2R4fSnNe/QcWnQ5UmuCA55vk7PSoI5mmY5G31WLh6zTzZ1+GYUc26On
PT4bdiouO0TPXP05oPzaInMbIag7mj3koKdkQZhEP9smUVoDPEP4l70yVdr7zjDJgf8vSUePI2zatwkGFeiP8NCVzrgH4wVT2nFuXRdGdDDURmYUPjRqNehFAOUhvM7m
sAPAQHqsHgYgHIUjqZ777HEBT9vsO5OYru9h38RPNfW02MgY8fmqdymGRGSVvkv7bymzngLMW6igjn+CMznec9IbrfL6baMuCl03bPAgR8Z/WBj66qHeFjTDlz7FArEt
he7Ru3PZfuvJn7ZlhGFd7oqsU3wP7y27rUvq012oXFKz+b8G/NvzFIFLgPJP0OMvaosjbChxdbNEQrZZIbFSZHl6yzhVLlcXtxiohkB0h/P2KWIx4ZzW+jXnebID2kmk
qHiPWn6RMDizHP//ZqweHoM0ksEN8pDdu1qYPp/C0o2wSoavkXA3OHZVG/s4ebCbHzK4r0hbcVKwJciYWbIlsiYpJYsN0pmyBFSqKQ78zbrSSu3pf3ffsET+Xp5Fotdr
pFOiDarTYEHmrP6vSYdqC2Ju4OJ43r/pgsYnaHd3zJKfjkzDkB17XP0lDom68b94KU2v33iOd7TvCMBPfY5cEkdlVDCQIyUXoYHE+YRIk6D65UYmZqLCmU55zJxOLlwu
7EXOGu/j8vMenfeI3AE0TtoNDDXqyph0ydP24hLnf1UBDOLOYkk912/6aCZnWg14qoqt1hHZxKQOdi4cOT2yU7gMuxsSGrwiqMSs6EZ9iU8ZiKcd6SH68mtiXiN1/Whq
4Fp6WJo74ahkX1EQe0WyzMYve0jvJq3tL+g8PcFB4EQaS1t24yH06NnxN5rCyLa6b9ViXTIYwXjJbxedLxXkZomAIUuUxwKH1vyj5FhLVkQBxO8XyDCigwqYoCu/mbTw
WTkEiaUf+jbkNOGegJf/2FCdcPjR5uCUFTJ9LC3i1oAJU7zlO//kzgDlkwfyAXj/BFh31V5Umb4eGuP9i7Z1evetSo46JNIh2FMgyDkdWK644yNWTdVx5YqPHXQscTC/
YUZtcAON7DwGC6t7LnfB1YSS4TjgfiV7flsDOft6DJtHZVQwkCMlF6GBxPmESJOgh2KtItKt9pLoSwM1Kj2itZoFbwkoCBVsYFtG3NaP2NeTD3zGo5CtQ2cCXcT2RuvP
5qS7Ib4qbJzi/RY6onxXdlCdcPjR5uCUFTJ9LC3i1oD387CV7IhZZqTM8jElr8fibymzngLMW6igjn+CMznec2Qj08d2PzSjY5kNB3C4/INQOev1S08uDUJEl8uHZDdY
qoqt1hHZxKQOdi4cOT2yU+HLzIzuDt/96ESLJELfIv0oiEqze0Wj6U3y8Ga4OvQFlWMCKy0RgodN2P/AcYXsjPOYF+5CcC0l98qNKSO8HhzrszJROkJ5xjpZtiXUB6rR
tLnh81K/zzYJfS22gUxKNGd01WW/4c7eHzRnYEarJtnxZT5qWXn/rMfxXMzoEkPxlShWgJzQUbnO5j2K35n2mGJu4OJ43r/pgsYnaHd3zJJjULoFZVG2phyu+RZn9qpc
uGMMYVmYPw38oSKjtJX7tIRwugVV5qoH09dInWio5zuMEx1Ue27/nT5d98pLx3k0AQzizmJJPddv+mgmZ1oNeHCn52qjiKgg2jwX3IkcxNjK6jrgYCuZPCvgmNcMFLqP
wp0PVoSth2KPEnSAsr5ZGSPYG29Spj7iGs4cxMG1MO6FHEjseXx6247STIxngcjXsv1riEA6t/lBrYNfoclCYHMP5PvdQS6d59Pi4fuJDR8tJKlWrRjS0ROg5VPxK/VW
i5mZGxOU5HKB/TD6NnH4w2Ndh+Cnj3o97Prcvsx+iXBnwPsQGZmV7OCeg7dhKXBNCkhZWYV7SGrnjv2J/n8sx72IzRh+00+UhVUC+yIgs7QOgBkDSbLk+rrCK/QQ35pU
he7Ru3PZfuvJn7ZlhGFd7h1QdDnHMlJwWZEczJj1HhWBgUFuNKojtj09vVZkkmYQIHxIkXCcs4QkXucv/k5bT1rpw7OWA/9/vt78DiCX3CfMa2oT0L1QH4oJO/QODcaP
BlokmHMShin2Rpqbu0gMx4ClZecV2XUp/p0C5+ZPWAOl157nUWNGXP+DQGYDXD6nCffOIBwaRBuG2NwxO1NLhzNINWUSh7QcKw1HDViXWal/yTpUl9lgU7cRPzQtMccd
sHnLa3fp7VfHUXI63xLw16+L4P6l8C1qwgludTx+13mZtEM5yIRFJrmZ96T45WzFNEUxI0uSUED8YFFSElM6A7u2SgjQah3pXA65VOI6aRbX5/CLRqVUhn2gkMi6+r5v
+2S22zXJLvkqELVgiKbGVlzZdrIKnQjARNWoxB1WCMUlfVEhCUuMueTF4nXnLoVtDZhX0piliffOoleE9EnYN4Wl2ikosWdUHCZstuksaWnLTTEgeAldX3KCBLDJ7ZTY
wnCr1gl00ecZ5/KOcDeL9lL+BVpuC4scikNlrF0z1rzP6viXC85LZHh9Kc179BxaAnLsVkKhVCF+a3Lri6YOm4GKXU6Kwui6XPYvhz0oQS+fXellLMWKE3M57P+YLtYl
gBwj73huZXibGQWvyZa0L/eutxu/ALL0enStnF1grX788TiR3idYp/M/Z2fR2hl4nPS6Ccvz8AR2Blj7NxFLJ+dUNNacSz7xf9D+N4c8p2MQI5EF21MS0A3jyhdqNlrK
30IathBidJFS99YPmbt7yIhh1+hHuwoFCqkzayXVhyCfTxhUnbYbm96cxAZjOtGUaKSWkT08c36ml6cbODDsZouAbcVumgfMm0lRxQdxnSSrRASrYu3d6ddVlgit7Kh2
KKDL9W8h/qWxTQJnRRrV1crlpgP4VUiHzc6aQStnEOZe7/rbkx4ke88CatVtzKlOfGefOhCNlWSn78Sgl/+cUKedwGUujgtpecUNsq8WJjku961vv60vs7xHPeT6UvU8
yuWmA/hVSIfNzppBK2cQ5pqigwoIkBBtp5+gbb+tp3R8Z586EI2VZKfvxKCX/5xQp53AZS6OC2l5xQ2yrxYmOTL3h9xlVHg5woogrjMC1SfK5aYD+FVIh83OmkErZxDm
ta7EBgYKGdytTj9tJcdQfoIRj66JR476hS69hiptybP2IVdqnM2Rwk6bc0xAW+VmQE1h+HIAlOeEGvfYXrovB1Aq4Uwy/nVfkTnstUHu8JtcNgfe2xIxW5816s8Yunrs
LrDME2sRAJu5CtYzIA1wiQbiPu+6I0jWW/AGObhrZ4NoYkzi1yOaOxGHQWGO5Zxsp42ATNn9RTash5bE39lhgydP8rT/tOhRno9DEoHffA9F5J8Hd2Q4+9lt2trsuGlW
YUsXtSqmVcTyn5/Ze79JM9+t3MBIiztwEUYRMldJQutTYJWxOfQz0djbVWNe0p+qAwmaz3cdTqI4NvHj0a/R5LLJ5EYfrDeJ3h3R+x82qtVn4DNiwpDuo2Fey4qyqTb/
MRNsrHJLsX5uYx+GyibWjs3OqvbosFkAM/spQ1QrRbLmdPwjxvfEZFqHPygryHua3vc9aqxMGeFpaENZyuJ9gNSOaIb+UFCFO+it5DgLXSf7rYOYzgVtfkRqqcU5jdlT
a45AQE+CvRbtELf1zPnpojNbotBH6tf3hZ6F4flblJFjHVakkbtYP8iLpG2slYx4IjE1GaB+QnvN5t/w7sK8yvfWVPSHeCpGI/o50UtVnKnFXsZZIzYcWW8jfy674uEW
wedYTg+t5Z83M+ce19jArkAQ5jbiwiRixlMvzCK8kkRba59b/oVzuDVYnVbbO+Nahb7NBUMJAj5WnkvUVcUuPQUg8mc0P4n+aOdBuWepQN9i2RIWkdaZQ830XyjwA3sq
+g8x76faacnRA1FeL0hYlDZdRNnLhs1TrUXxQv6suIH31lT0h3gqRiP6OdFLVZyplgasXs+iuxM0U0WuotqsM7RqHduNBYNLr/jm3OV6nsNAEOY24sIkYsZTL8wivJJE
I/jooot0bvq+VVQM49CuIKgPeRSiiiBSLrNM6L/oJvYqvyi7JE/ACnuqFsDsfZQe6yn4Ac0ibG7qLYWTTOs7htsQws340GaeJMAHLzfWw/Vh1PpizIHCvbB3w691ahiP
8aueeDpm6fRHb1mn2YrYv7w/4/fsFyhKZLrZnhI5VtuLJ2V2PvCiEGEO+KqrUptQ51nvAjVdF8k5nRJzW9yKIQ2gsUZ+ctqxBxL/aTMmaotTz0sQXH3MVbtV3cZz0HlK
i5msU7Df7NxAcc25o4f79TkJ/s9u7Gk7H+f7wRicrMZVM0nDvPiBpGaZRttBoTYtS8EgEux70A7NVBs/T4hvzNILvtLImYKbqdQNjKCXwWXW0/BuHSseypfbystP460n
3Fsmc2Ozh3tLaz0UxD3sHzFVeOElCFC1hNfQ1Fqu1ymQn+2/5fe7PJMJvVb5UryRrqOeo4ZWDeA39MOVfY5CJ3PzkoY4J2AwZxy4yEkdqpH9gCA/Izj6ngovhUkdq6DL
yOZWpuFL37KAKDjFKRlIlBCJLOS+HkbD+vejgUAUYcESJHaANvR3/LgKNPs9OH+K/AY6EnFsaW4kH+LFY0z/i4jmgBixwWC0DlkXdJP5gxYdDzvCjNT77i2NpjkAPOm8
3LfhCJrXLiVSzFA+Vz7hwKlbujJ2gQjMrLlvPmxd9rSQl7R1G73J1Kx0A556GbKOCmZOSH0xeWpvrmnBHi0qHaL+8sBAYnDeYAF5dFVjshJMMG+S+OqSgQB4RI4XqgJG
40/zbOQy3dj9WAK3fmRLp5NodfSYJSB5REA+yq3lMq7e0gekjBPQlP2V6b/AJA00UOFJwZAyKwEwZu7HtI6lfCLLwxMrtW9oDHpbiHkif2ZjaOBfRHyqNuMrSu9KVCHY
y00CmsMoVk6tKs0GddplG8P1ukga0hhm+DOEydkp28IVqfC6IKN5VUD9pyVi50Phx7/4b2NCIuZEKeOqcNz3o3cKHOea/3oW2mxojccDIZRPpn9l5Aw4aC52FIsRpNYK
GAAhuM2Ni9ofyDfTayGPLrc9nJugUDyQ/GtmLbThYwc5Cf7PbuxpOx/n+8EYnKzG9Zn3EjDc9IdlzKc19l7P/y0prabbN8zBdagKQBdOqz3Nzqr26LBZADP7KUNUK0Wy
XbAmceryv/eoD6rA8WpOwjhdotvHM3Hl8PcGloeIc7UTYRTXIPmMPCT0zmJE7MSoK3Q9FI74kzvLpodIK/emJetrHVCQRpp8CAK4u893V2NmMajDeAQLJlfQVfXpQO9R
b2c/FhwgFm76cayrLhJAP5cPjm0PBrMq0IQjBn5Jqwamp9epKmGNBRmlJmMfjKB9iydldj7wohBhDviqq1KbUOnHjD7AWFHSApuHjr8L7MZk58NvRg5mXKM7i7uZVmc2
8mr+y5OntyBQAjLdeJoeLjWtK0QjyrszZXlu8AdYrqeZOMOn5JyLetyERCpgFWqB+49DwRDJNj/L/Ros8TL5BbhXCLQDLm5KOQNz43YlM+meYWjzdzwhrNDFY1tx3p28
CnT4yvPoQrqAtWAmfLDalk+mf2XkDDhoLnYUixGk1goYACG4zY2L2h/IN9NrIY8uXEND//qkHPWZZdAlEp4S8rRqHduNBYNLr/jm3OV6nsOpSftmmCtiRG8XHNpLt8uB
m9gTYeeU0JPm/IMCBezRafKHCLJb8n4win889g9m4l4zvoMGCmapTBhPqcx+SMtpHQ87wozU++4tjaY5ADzpvJu2800BeSzWnl/4Nt0ott2b2BNh55TQk+b8gwIF7NFp
McDcrS/rGEq01gip2YmxVr1kVCqlYRYZC07/5l5IFE4rRQPV9SFNuPBfOqrVkV3mKau3PQ64zW37J9ZqH2zBUMqIJtEmvYeBjKtfeWMCbYhvEzpMRx2mq75FbMsTWyTL
A6EvQWzZXRgKAFppQ7PQTjlrf2hXCVN1zEJbu2INdUzsu+XRgGdYrulj7mbX0+Y/3tg36JZIjTN8D7VQ9R/VsovzsVukaGa6N1yH+UEpqbUeZwTMC0/rBJXC5QKs6vNw
ZVtNWlDjWITAoKtmOqXCfD88888RZUDAVhXohezktK+YzIYE1Bdj+o6IxcC+awzdDyTFZE+koBq1JVGxGMCzPz88888RZUDAVhXohezktK9bQcEdbtD9TroyKie4PpYq
4/25HNQScdN4m5aLMSJBTKH9khJ1Ld+9SrO2jJxyM6a19CjabrqRMro9cdNFJqzI89c1r7FRoQxMnpH67y0P40+KPsnBYzS2ovnuXxWVg88J692gkwUnj5b0rLLzhEo7
7ABd9NLZo8iPi9pOOOECdmRJJY4rk7InR/dwo4V7KRAxYmf9TfvieZq4i1+4laBeWbdlIT08jZtV5+9pALGQeYtoT51Ej+DEPL+tMJF4wiahEPvXK89Tua+1Tqgiathh
Wazflag//GrTi+1JwdCAVsRZREfD4DCRAxyoLEFl05KnCwpeuiCDLqLb76DEbV7A5yH7G10FFC1zNWcVIDN0k+zkXKXgYPEtXBbwR2bKIZy+J3u9Z6576Fh/2BhZlyMK
CT7ZyYGX15Jw3TY73d3MECKRPmbp+4ZenCXHPSTu3tX3WC4VuzxOuaFcTzLTt8BnkyjNbvtloOMTsWlhkUC+Sk8Woa3vCUibEu9EBQGxg62ii6bAVrvDv2smY3SbaEo1
2/kCIcUfW+/KLSRTCF06Y7DPrCzgt8ho6MTxoAaPvYl0OhPab6pz5K+2hX4yK+yZlwjP6DwnImBmnpEZudTVbRsRbg+GAwLq/HFndivTi2LAa8LG1RH5K6YLHhV04v4y
cndbJeS3PIuqsc3cSX9GGZcbJgrK8gqtte4y63U3BYFt2zIoNjgIt2HZYFeGgwEOfc0pvKfV87iSH5M/kT03ub0KuIatxtp8NrhtOQ7htgVLUjr3iuoXULL1B5RYD11d
sTOc571I6b5Dwa7yOErq+WSbineILPWvRlxeEBgbCjZBYGqn94z1JbM9nrhRSd6pqIj/71r3FoPy/gFoX56wNwugOaqV+M2g/WMz96JjDtJyd1sl5Lc8i6qxzdxJf0YZ
iYI1RWqT4bbdhd6bSfo7VmnC2llXrj9tJGD8TDeV74izrQ6rdtIAjDaNcBxTnr2Vi8AFBoHz9ahMckTWJlvAPtYktEUR6+2QJWBl2C/uZcvRC9sHbzS/0zlckMrn1MwO
VgYNqtgImawCHsNKfI8taYg8pD4HtnlFt0cTAW0fMwYJPtnJgZfXknDdNjvd3cwQIuB/07MIQyWMhqcb95ufYO3W5iufZM6wN+8aIXbsxUpEq1C1+b7qMK8et+yzMDA7
juR+xMHz0DBKjvSMagaI/EbQClGMsJ3g+BoXMRtM1e7j+ebu/uJ49LrADT3VvUVjwwF/Mln4m3pCt80+qdAEYvsQUBgCQV5UQ8qOjGTWSih+F2WbBE7feAWs2M/hij4C
lzAg3NuTojdT4wGlMX3Dm4N/qRvhWwjvKE0755rKsOtae+E4ZvabNXjS5z5k9hPlv+7+n1uFONHDClOM3nrtduch+xtdBRQtczVnFSAzdJM3z95avBRPyjaSTkJMg5jb
jitMcO6s3J+9TcMmEYXYvktSOveK6hdQsvUHlFgPXV0KOp7bs8Jy9SE2sLt5cE6GGmjeljmMnJqeThSwWIB/c97YN+iWSI0zfA+1UPUf1bLKDPCXgOaxzteBILbK9AaT
pKzo8TF1jr4G1BoKtRb9p97YN+iWSI0zfA+1UPUf1bLKDPCXgOaxzteBILbK9AaTumfcrKIXNsuMm3K+5kq4QYuSKXRQnA/hVU287DW/ftmwjdCGxT0NrIYAdhynzpfX
G3OfIDhGeUjhHEg9AYARbichNs4BkN0jWS/1+zhfKDyrUwG8Yx5ZsqSriNY3qvB0wIgZwLJjzLxFZV9k7f1gr1jcbbqhKyj4cSXVzmag5DAnPUyPFVX8cKpO+ySb+a3I
ygzwl4Dmsc7XgSC2yvQGk1+jO2C5jrCgWy8MvQxKvELKiCbRJr2HgYyrX3ljAm2IMrLiQXrmF47BvD8bv0Qq6i8gBZy0K0A4W70t/pya2tJ/FwudDKXKnFmdEuYD3eGw
rvq72+42b0UAn0s71XnRdMqIJtEmvYeBjKtfeWMCbYgDOawVLTVsvapw7M1SmG9+funZiqE9xG5L78dUkAocIcqIJtEmvYeBjKtfeWMCbYgDOawVLTVsvapw7M1SmG9+
6WEnLBIXrKzwBXk7qIH21pZH4laLr7JJX4Dskf328h4DOawVLTVsvapw7M1SmG9+smCI8UXnqMRhmfOAoGI4KWKRUiysamR7h4papXHEmjFke4lnB0Xu4uXNihjiU2WK
spxPSslh0PlZcZUgLjKU1IoGUojD6R6kD6uzUEnHGd3riIB2JibbNLuiEw9hIp84vST+cWS0Z7XA3ylj3MfTs67IJwfc0o2Lng6NZiBdODl0hYbo8KKSOp1yLqvUfql6
Q0AkG/TABuFBPYZEIyDiD5B/keYmgETpbFXygYEtO2pXV+7Gg+bU+m7D50AnaMd3Jp13af4CzRD8mAodBoynpeIePStPGhnptG5vwBOv6+bSJfOaTDzDP3o3UyK+yyXH
kN1PatxQLn6ARD8GGEf79cYm+r9p4OudgijCjn3FpKje2DfolkiNM3wPtVD1H9WyqlutNZcVVQzUOPxk5eMeBc3OqvbosFkAM/spQ1QrRbLJuf/Xv4LtLJIPNeBNxIA6
4h49K08aGem0bm/AE6/r5uMzaj4gad6z9SWHS024+99p9x/TVikdNR+F1KSEHESYMYT3+SAG6MD0oHdaA1+z7721jSWOnkx+HKg0SkmdrkDShsqnWU+UwZdOc7BZw8C5
EOc2TQhxB1ZJtxGACP3JeDFiZ/1N++J5mriLX7iVoF4Tm8Tu6eeH2TzAIvregOPAlzAg3NuTojdT4wGlMX3Dm3Ml/QcigG+SxjraxpZtiKdkGVK3EwlqYnG2+qloAnE2
exYykexcQMsrmn4l5cPlCuNKu+vRr9iY/1c+jmUWgC5W47D3lJA7/VDt8o9h9AucOKRTIcoOQCjYXL+PbmvuTjMZOhC5TGC9AHBfw5v6feb6IhR6hy1I7VIYb6ngJjqN
iba4RubG3DcfCeEH4bmUKtFigt/vqHtZccmL3YdKA2NoFEpadPMgRobL3I77VWBaLT044KEK9NWiFRvqZTlwx2OrnO9WuOFv6fDwnwaaRidizBcAYtI+hrXGaLBh59uh
QtkmfEUtH7Tn7bAuZn2X+9t5x0JfjfMFDltzAO/oYBAbEW4PhgMC6vxxZ3Yr04tiwGvCxtUR+SumCx4VdOL+Mlr/0J70Fr+atAAf+GGXDZJSibb1Z/giBPe0UMoruFZc
ixe37J3YHsqhFgvEbGB1c+3ieNkVkDS19BgQrV/O14CcgkNt5nXJtbSETGN3ObEtR2xPEdIx7xRpEQD2z8jxgW+LVzeAI4Yo6C+uDYEteq1PDA7oub98bVjvgG+0+nMP
B9msefxLXvUtIHVBlRVBMQpnjpc0v7qVkfGItH7fb925jnP9SIdSrCwe+Y6uV6lEmvMxzXJd41nwo7ygdzJ5tmnC2llXrj9tJGD8TDeV74izrQ6rdtIAjDaNcBxTnr2V
XWo7IirNrPezl+Y4cZL/k3sWMpHsXEDLK5p+JeXD5QrjSrvr0a/YmP9XPo5lFoAuVuOw95SQO/1Q7fKPYfQLnHWLGz1j4rHuTqhiyXlGFaaP5vgk8itbiF1FMhbnHJie
TE2LdOmo2nE974iJyIl7kuzGsXoNNrxFJ1oqSjVVaqUpoCcjQLwgXx5AdDZi55ce0SFG+dzIzIqeoUDYU9Y+n1EN0XFVS7qPH/APwydBTrENmrZDyi0xF3S02W/aDjdv
0e0TCPtI4oau2iIWQ/tOvrSi42CibOM+/jEPGNo3WyPPpFTc40rr6Re137up3YmWUom29Wf4IgT3tFDKK7hWXLMZz5ULbCOlbZsFhAwb+PldajsiKs2s97OX5jhxkv+T
exYykexcQMsrmn4l5cPlCjrVyWeACVZSJK5htMUy/x5HbE8R0jHvFGkRAPbPyPGBo2FwLUmHRIs29LcLivYgQCpB02C2d3hVYEehXKvG/KysWabwR5EwNHFY2u9rSWmZ
NBlX0T0Fb12NVKzc3NXgijiRfgujThAl2To+k00THY3dDxOLItr8uVdUPS31nd2RM2lbwi7q6ZAxuOkVWp1N+OZ2jxLmc4QF0IPRWrLsvXoZuQnm8lFv9aCY+kuktcmC
anQmLMGGUAUw6anMFwb1kMJ9nN8cgjno9McXhXRzuVtl4Wco4VodMBnD557HQylFiYI1RWqT4bbdhd6bSfo7VkLDPyK4JR7imho4e9Kk/3i+Lv86f2jIYwvHFdwcXzoG
LbsXMXnSslIa19oP6GMxMrRTkZtC48scT3y5SOBTyi2+tQ/TWMTO0g08Ye7CQuupiuJ4DiPrubHgEpeMHkmwouaYMjAvIiqWqE4v7aV7CMzGMjQppLQ0XTtfm6oG7z1r
2nwprEjEJ/BEkk9longSKcqIJtEmvYeBjKtfeWMCbYg2RdNBn8k4oZiZIp0xLMP/yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFG
dQAftNleQV3YzJYHykVbBzLhxmhYqgtFWuNBznYYskuaoyxNU8fuOlDDfHDLcZkTQWBqp/eM9SWzPZ64UUneqfcMVb9Du2tn9PvPwFFFRQLKiCbRJr2HgYyrX3ljAm2I
QMmqsJAIM6uAKSZME0akDK4tSJoZJtG8yI7ZjmwIBI3XJ4ps8BDtBhJsiekfumSSFOAnLeaNF/Ymkft7tZkWAD2r8LBQWL+vmb1AcQADKhPKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YU1K76Ha/tLSgr2aD3/B2ZjPW8nmRS1gc+TIjnbkupKBTBdsaRQTyE4hC+P269u1KXJkTx38zJquLieRZiUlINh
3tg36JZIjTN8D7VQ9R/VstMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o5yH7G10FFC1zNWcVIDN0k8LyT3RKeBcg+5fDaYawF8SZZS/uqXK1cW2h5KwDu8k5
YAyEzu4aubwXNbGVPKkCDMqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFGE4mP5yBy1Ghu54UO40JYId87eGsX6gYkvacBj9HvdZEdv+6giUNSzAdHJ4f+jWFY
DGGjYSX/mJhUZdMFPwZj1uWP7lDFt2H4il24PqGpNyrKiCbRJr2HgYyrX3ljAm2I9rswH5Rl3UkeJz+f63rT764tSJoZJtG8yI7ZjmwIBI0qcgwH0px9kdX5aYCIw4ZB
FOAnLeaNF/Ymkft7tZkWALYMzw/JelQOwKYe0PdIp+MrcoKAYE/dklAtCtcR7Jvayogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YU1K76Ha/tLSgr2aD3/B2Zj
pMdkvg4aePZ6Z0eyzw0cIjBdsaRQTyE4hC+P269u1KXOH2FHC2/36yb+3GxaJayplmJwqSxzcxgAuF0utn7RHtMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o
5yH7G10FFC1zNWcVIDN0k65ehsxIxa06CYZd1n8TBfeZZS/uqXK1cW2h5KwDu8k5NQ7CUaYabiy76FywKNQdrMqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFG
E4mP5yBy1Ghu54UO40JYIV0l6dsEE6OGC92mx4JraisevAeDKZ5zE9yFfUzDVIYoDGGjYSX/mJhUZdMFPwZj1tmz6DqX3E8GxW9BW62gmorKiCbRJr2HgYyrX3ljAm2I
9rswH5Rl3UkeJz+f63rT7704fmZioao2ROAG4nqc8V7KiCbRJr2HgYyrX3ljAm2IaS0Esno3/wPkQvGBBF+bZacLCl66IIMuotvvoMRtXsDafCmsSMQn8ESST2WieBIp
yogm0Sa9h4GMq195YwJtiBJGqJWn1t/qGroimMFAGFaS81QA1hhc2M8LHezDl9Kgyogm0Sa9h4GMq195YwJtiGM8xTZacX2EykrBdtIBYYTKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiNMhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbgMuiA/7HTrnioebM8Y4bRjsqIJtEmvYeBjKtfeWMCbYgWMUz89adlGFsHu89hAjcH
7ABd9NLZo8iPi9pOOOECdtcnimzwEO0GEmyJ6R+6ZJKhjhkW0xZR4jr1EKYyTILNqJI7YEbeIAYkNBFAqjXCBJcwINzbk6I3U+MBpTF9w5vg5F9Xv/IMzo1gV8k3YZwc
QWBqp/eM9SWzPZ64UUneqZVYURojG2peArvAJeQcrWw9byeZFLWBz5MiOduS6koFQMmqsJAIM6uAKSZME0akDNScD1CgcTMtq9SDZI3h6qOxkdubgOAyfgyIxZC5MrTF
ziNmgl6L9delvhB/43lacacLCl66IIMuotvvoMRtXsDnIfsbXQUULXM1ZxUgM3STwvJPdEp4FyD7l8NphrAXxBJGqJWn1t/qGroimMFAGFbtC2jidYycQaEjacfnw8oE
3BYAA3Nu0BMXtZ60286uGtUSd9vOFccXpaTrC2SBvNWLaE+dRI/gxDy/rTCReMIm3zt4axfqBiS9pwGP0e91kXQwlOUavYDeZsZAsAOQL4iSNw09cGng8UC0zuarcnzV
AsQvV7RWFsAF1HP9qG4TMVumPsevnc/8arRqisxmpH0WMUz89adlGFsHu89hAjcH7ABd9NLZo8iPi9pOOOECdipyDAfSnH2R1flpgIjDhkHvdozjhgvmPYEbZMFRW4kH
qJI7YEbeIAYkNBFAqjXCBJcwINzbk6I3U+MBpTF9w5t7Nuzc6TRyG2pDcU4UDg2QQWBqp/eM9SWzPZ64UUneqZVYURojG2peArvAJeQcrWxcb8eomncCm7feOC1DLKVx
QMmqsJAIM6uAKSZME0akDNScD1CgcTMtq9SDZI3h6qOqkPVAKxmPIrVeYUUUWch/aS0Esno3/wPkQvGBBF+bZacLCl66IIMuotvvoMRtXsDnIfsbXQUULXM1ZxUgM3ST
I8XZSVq+8r3SwyDHpQhuOhJGqJWn1t/qGroimMFAGFbtC2jidYycQaEjacfnw8oEBoytnJAlkhAUaJHvWi/jRtUSd9vOFccXpaTrC2SBvNWLaE+dRI/gxDy/rTCReMIm
XSXp2wQTo4YL3abHgmtqK7obXfpHW4QxkfrxdN9Afp+SNw09cGng8UC0zuarcnzVWAkV2JcHjGJZwDKnjqpgf8qIJtEmvYeBjKtfeWMCbYgWMUz89adlGFsHu89hAjcH
rkKKqZIxJKZEJCKIRWMNrMqIJtEmvYeBjKtfeWMCbYihjhkW0xZR4jr1EKYyTILNUwmRoUqzOeW2UvYBJntSMXI73gMzvv+1OfGMEuyVGhdS05M7s90EhofheSI9h88a
qxVBtbhWvXS8QxWoBC/M18qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I9rswH5Rl3UkeJz+f63rT79VSeWw0dbitdHCRjL/CYqMkVri564ZJXY4B+X0pLt2Q
aS0Esno3/wPkQvGBBF+bZb/u/p9bhTjRwwpTjN567XYM28K55L888CVmb0+UBGteyogm0Sa9h4GMq195YwJtiBJGqJWn1t/qGroimMFAGFaL9Cc7PyDE4nqTgZjDyP6Q
yhv2DAx6htG2rwiEmWl+ZdUSd9vOFccXpaTrC2SBvNXjIW+L6/aZ/r4KuyW5BY9U+/6wHJX7oql7hVkSDDfsfPeejjX5LVfeAaZ/Z40rzhWSNw09cGng8UC0zuarcnzV
Cjqe27PCcvUhNrC7eXBOhjSXFZ5fJwtpSZ2s2O47T9kWMUz89adlGFsHu89hAjcHDYNsnSXTYY5S3BjV1BTk5YCmNxzirTYd7fXcs4sXVIShjhkW0xZR4jr1EKYyTILN
Nju9CP+n7rhpBkS2pegxjpcwINzbk6I3U+MBpTF9w5suEY+SCWQtHS8LroBVDu2cQWBqp/eM9SWzPZ64UUneqXFa/2wetEa233/PD2aFmReQg+6gIQByB0NisUB8a0Gn
lzGVf1g75zdPHELQsMdkbtVSeWw0dbitdHCRjL/CYqPj+ebu/uJ49LrADT3VvUVjm3XCxw5J6ro0B8HbB+AleL/u/p9bhTjRwwpTjN567XbnIfsbXQUULXM1ZxUgM3ST
C+I1SZr8COPCkSQzuNQcZxJGqJWn1t/qGroimMFAGFaL9Cc7PyDE4nqTgZjDyP6QRHl8A6pExkjxxo3VttEVldUSd9vOFccXpaTrC2SBvNXjIW+L6/aZ/r4KuyW5BY9U
uTw6wpEMTT1pyef2HB5y3sYrrLBxLv2TQGxj8BkGeNKSNw09cGng8UC0zuarcnzVCjqe27PCcvUhNrC7eXBOhvLPckPxCsTkVJKWJkhhdI4WMUz89adlGFsHu89hAjcH
DYNsnSXTYY5S3BjV1BTk5Sln1+L6a5jhrvLK29hmxHzrePAePgZNPRYPYWBd+Q6iNju9CP+n7rhpBkS2pegxjpcwINzbk6I3U+MBpTF9w5vxcx69sXHprtiS4fE6FYZ5
QWBqp/eM9SWzPZ64UUneqXFa/2wetEa233/PD2aFmRfSQ43EBgKroxSYDs3ORJtMQMmqsJAIM6uAKSZME0akDNDPY81AOZnvZcQtLD1UDzHKiCbRJr2HgYyrX3ljAm2I
7M2pfsVdKJjxQaYnzkufkAnAb4QkreZc8z0CyBkNBKbKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiDEdVthgIYrtPa+D4s24DDyAo79L2BhBoQd4X80WK8R1
yogm0Sa9h4GMq195YwJtiMRG1849/TeWFNleaMtqMMW+Rgtf+aIwriJGmjgpJ6RXyogm0Sa9h4GMq195YwJtiDRYlTE78nku/iN2dKkUNF+EKi/qBiGRTIbY5OBnxaf7
7LJUgQn+/UTuHmCHZfw9gG98z2RRPfwkjyMvxxcG9oBakayZvZQeWDKHMzNNrK2a51KgN9fIe46DblhHF9u30m0ILZFy30U+pWt6XvbkSahAiKaq7UmP6wJpP5JCmOLK
yogm0Sa9h4GMq195YwJtiDoLLRXFdl6eoHGRGUt7b0rj+PkMZgKZDmvR7ccXURbDbQgtkXLfRT6la3pe9uRJqG041bPemCZq7oMhKVUsZMRw70Un1Q9IUc6G91GseXXA
6HcqaiYxO3xdTuvKeUVmXrZfejunzBU7kz5skaK+D3OWlHJXiQ7Uktr2AI42n+P1AYi4GCI3Bk712//+HFVPj8qIJtEmvYeBjKtfeWMCbYg6Cy0VxXZenqBxkRlLe29K
rmBsLlQqbsnR1McDETxFqZhKrjetMFaGwe1a7Me0rAGNZU3zfLjTNGmBXIKdpg6dyogm0Sa9h4GMq195YwJtiDoLLRXFdl6eoHGRGUt7b0qkvHD8y0IY1z49L0JReCky
bQgtkXLfRT6la3pe9uRJqJuP5XOt9A/iBV/NAZvdP3mLYGtvY/Vs1h2pytLRB97E6HcqaiYxO3xdTuvKeUVmXt7OSLHo/yPjCMBYS6NKboU437pqpXXAAj6jui12kHWF
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYg6Cy0VxXZenqBxkRlLe29K+3WroLhD+2OPkb/8JlBOhNix8eE/cWgfN9nJGUtscdQ3u1V6Iuk1Z7r3idSlvT0D
r0cGXd1XYajNa8l/fJ5M/+h3KmomMTt8XU7rynlFZl7K7FdidI67mGcGTR5s2HKtDNZ0GOC2J81lXrvX0AbZ2Te7VXoi6TVnuveJ1KW9PQNXtdTnLGoLlVMZpppn1bQw
PJ1TdigyexGYeExcgbAzzKfj0tNflfIY2g3vVQHPdT8/+30HktiLeje8OFfSG0WJyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYiYmKLq+tHjCBCvnTtS1ZNg
RFue1lt5WoyWIkbZNEwcfG0ILZFy30U+pWt6XvbkSahWiw9Y+cJNNb67y1nOzzZo3GpZ239z4KDh4Hnpd9UBXGYkmqYAhQ/hrupzHivVUvoGgyIc/DkbJJinnUgBuzjB
eoo5qe0z7B5PK3RvN/DS+k2s57Q86Wae8QfMbcO4Bz7KiCbRJr2HgYyrX3ljAm2IqgaPkw3YWtsNAYYfrF10SzdznC5JYvRTd9b553cnJVbsxwgGchMz8VS3j17TJtfP
yfD4Ai82Av1anYKXUvVrL8qIJtEmvYeBjKtfeWMCbYiSgbT1h/uOSGcsotORpa4A138JmrxVKRKGUH2AsswEuqXjDm9LNiX+nxs5p/yygbeX6IwZnvP00qPbTAgjhr+W
3qryrb1v3B2w2k0mRwBxBu1kZn8UwSFaPkMSTtF3IQTi/zoSeMRAlrGxUZbCyQl3YaBeb/oSptenUn7nWZzKIMSI7Bu0pmrXLZDwBi7Vpq/a8gk0x+3pzHrDUtVgrbbc
pPxYt0hZr7GEUyg91r6vpVlCD5X3643xa2dMWTzKqJ1tYl4wH1oGiBPPr+Rxty3EQ+w01OJJfKh1N5LQB6682Au3Xq2kKv6D7XlRulaz4k8A4PJir8rj0cDesxE+Ubt9
ALUUJv57EeErgSrG8iiwms0tWuONOKZGTPPdpRHyekpKnxyyElTNAM+c0BRAgdO6tDAWEGu73936EVqbQ/LXBoFIw2MZsfxVs+uw4O5kLyQtXCwl3z94rKBpv+jbDmpP
3HiiqxORGxM3c59XuWKDmh6vN4Lq0U22nop3r92aURwacmEEXl0nYZCwdicY30opAzmsFS01bL2qcOzNUphvfirt6kELSYuU45P5N4tFqV40MkLmFYyJXZfglVK4Cw6p
w407nRthPzi5jNiBVln7XFO/vCx9Q0SxMxEJVGttLb+w6cUXOTrd/AbJTnnPpsO5xCJZSSNX65+OWCHp4QSkzXGt84nU3fwzhDtkTDJttxxATxc8SNKtxrbmyGQ6aRLu
BOdO8YI+T3Tn9v/MU6z8zKXF+OQveKBzy5CULZ9WQnREYFXfdmBKHj+n9KamUGttg0Lwv5HdHDYSi8iXxf+DHalRFYilDzJ7TInlYsiVdR5NxmPWZUBKgtKuE3hcRxzs
gQ0pUEzetfjxrXJrsqudqBgYwKnSMMtuEqUmXYi7DNEicoDzFWo21WSc46CjTN1+5xNVsfcv/eXvMcEWcz1GB9ryCTTH7enMesNS1WCtttyhq5fN9GjS+Z8p/vUrT4po
LOyFES+eE5x9Z2sGvK5MWv9SDCuTEG2CfCkEMDGRa2CwSoavkXA3OHZVG/s4ebCbhlD0yJNQM6ZDBejqGRP7KYNC8L+R3Rw2EovIl8X/gx3uh36zywM2kChUQ5hH4WIB
NBFUtuv9JvUuOuwpUcF/5OEVeYBtHot7eYFbO3lBiAGl4w5vSzYl/p8bOaf8soG3nbpec4YL13zkLQZRpHsg+IoV1OeeCXlNOM0cLnRIKA38HB0WkRZGrtS9qT9h1Vpz
/ArxS/Z166l2bwIqCG9P+1dX7saD5tT6bsPnQCdox3fjeJ6dS2dCt5GYSZSt+EBC12NmXCQS6YVNApU9GI9SAGNQugVlUbamHK75Fmf2qlzHl/wSRXGAMwbFJf1XdWi/
iFPPD4QgoGvDokhiuRnw6Uit/PondToUcWdBkmKNyWDZM6/UfUkOBx1CLFP+gdDDf0M0Q2r+Zj6jwUpVp1fk6Z9NVG8xFYX+EqTkw9Rr4PiJu5L2dzvy2mt7AZCfvsjW
SgEQuSBNhFMpCWNGJR8ChSZX3ZHtymEDth4AEXEolqOPkcrqb1MvZg/82Xc6BG1z/BQdtRhNegvPf5WZ/8Zk3uCj6NJVi4944zLBEJow0+RlLhPnjDDBFwR8HUwhn6K4
9PusDK/R31L38aZ2Y5hOc6PssD0mvrlD9BSu+8GzgIMpdiysd3WwiS1ttAFuPENZSSxaF07Z3lMEWvWuHVa9K+SRHZ+Hu2wUSu5F3uyuI4aIa4gwrDgTJdOv6S+vY/tk
QWBqp/eM9SWzPZ64UUneqd6lG7JFgUpS/JPCeWAYcKCetK5lpYpwfP0PlYPRFTYuKeTfmmlJfMu9W4YD9bRL9YFFX1TlakxZivDqOtSJuTSOC88ABZf9UzRlnaUbdHUX
5PEMVc0V7JP60ZlyyHKrf9V/zDEhi8kSWVog7dkNHVG19CjabrqRMro9cdNFJqzIaVnx9So7NF/Lp3rxbR1yUrPwMN9wRAMX8Xv7A8KHFS2XUdrw1pouU9icDyi75rQ6
+J4wzL/hcfXsK+z310otLpWlUrHciYtell3CmWzYIndlpgklHE9sH251GPP/pDBvYqC0Gel7V/6oM1+f9dK3K+qegXDySlr28Jpyac0ZaXY1vasLx02PCo6rdVBZiutF
V4tl9+TngaCAIcMOOSDydqfsbYvX6AGXwWfk3BbwyNrK9estFyUhZMvyj57JLqKZFjtsiWbDlUAEGSjGRfgZ8YuvJlAWWy4O7A8/91HQb8JMxH8N0qYu5HDwxINrWM23
v5lvBiZ/+BuedZXODZO54fv+sByV+6Kpe4VZEgw37HxQyyCtK4KKo16lxQoMAKhQlxsmCsryCq217jLrdTcFgWnC2llXrj9tJGD8TDeV74g92i21UoCf/2mRSzUaH6OS
j0ZpTubWtf85/NRNt38frk6+zkmvG/081Ok29a/q1gTp+K3gLrfvtU67bRoPB4QvP9qrET6eF7PH4vosV2V1J8MBUSLi3Sc6sR7Ti6N7EWc+CWQqquEZ9iSQXtlurvt6
5yH7G10FFC1zNWcVIDN0kwYvYgV8Rp3Nccb4UOlHYwhLUjr3iuoXULL1B5RYD11dAsQvV7RWFsAF1HP9qG4TMSOKq1s4PQ/dNxM2Km3rkh+/mW8GJn/4G551lc4Nk7nh
BtVChoKqkjuy1B8XJ3mBCqNsPhPoDqQ39JmpturJClSXGyYKyvIKrbXuMut1NwWB3FwpB767aQ0GHP8+04s+2ujv19m4lQzlcdDKNReY9oKPRmlO5ta1/zn81E23fx+u
q6JoSs8TSAc5Rds/X/Oj9wk+2cmBl9eScN02O93dzBAikT5m6fuGXpwlxz0k7t7VfrkTXLQaQ6Vmsy/zt7vH+b+ZbwYmf/gbnnWVzg2TueEqa15Kd4aC90Md2ZBvB9KA
tF4rNi0atjfVllKPiqNNx5cIz+g8JyJgZp6RGbnU1W0bEW4PhgMC6vxxZ3Yr04tipbcAlNH7GnXJVYYN9ArqnYl3YNcqp1dfw6l5rgQXh648KUCMaJOezbOpAOVOSBnI
QWBqp/eM9SWzPZ64UUneqZVYURojG2peArvAJeQcrWxBZ5adaALPCoktafDAgfIwSDdlM+j8YNvoYLZObteNbH6MSJoiO9KYjt4cz8DMwEI8ARkEyw93QWc4NlAtt24E
vxlnUZQTQdaZH3sh4+EurKCgyYak195MiB+M2paTxIfdFgeZ90EukbxkFYb/aVvvC+ejDj2nSA+VQLVH+ZX9afieMMy/4XH17Cvs99dKLS6VpVKx3ImLXpZdwpls2CJ3
ZaYJJRxPbB9udRjz/6Qwb4hitSiIFCP9+QxE3OI0Y52pwiMd8w2US7eoqibI/z+xRRHPLWbYozHaqLUqktEbzmv7GbsmFx1fOQioGcKliIfMrD3VlyF325zE7mZMXEcd
DZq2Q8otMRd0tNlv2g43b3H16ffqSDxA+9gDPQKQCr2/7v6fW4U40cMKU4zeeu12ZpwoGpA1+hS+qLxJLyHm91licIWaI8bjUl1gDr5+xF1Sibb1Z/giBPe0UMoruFZc
hJabJZBmEoLu+8liQRqDYL/u/p9bhTjRwwpTjN567XbnIfsbXQUULXM1ZxUgM3STBicAJpy7fPeV1bA1I3vaUw2atkPKLTEXdLTZb9oON2+xkdubgOAyfgyIxZC5MrTF
CYJdjWEovqN1ETfg8/TTnVXEycSPQmfVxM4FhinMNFdxEdMH3nVWr5ur4JTq9HjMw5533+UdmXU79TTuAIIPkB3kU1lnlKtVMD3eYawnIH8hPZuYVpydltCmziaeDv5D
6fit4C6377VOu20aDweEL0Tb0PckcayTEhQPYxa4EfAK8AiKI29mzCpW7jADuviwsYEWCpiKZFmyt/m1rByhGol3YNcqp1dfw6l5rgQXh67OG+h4RVolfTf8t26b72E1
SAMFWEXRp1ExlbkULe9wx7ubORLeiDWDVQfwFIsRd8TKUKmFmE4ykV3QpSzQenfjaek5tt3ZtQ/+hNykPFPOnCsv78eLjGPJjPHZxpsB2yilpjXeIAy5gaEepyEkJMFi
4yFvi+v2mf6+CrsluQWPVLk8OsKRDE09acnn9hwect59Of0PtwdU4UljFNEAkYepexYykexcQMsrmn4l5cPlCm84DEQfELwEMHpsnBdZRftIAwVYRdGnUTGVuRQt73DH
u5s5Et6INYNVB/AUixF3xKwyzAOh+UKBrTQSgRtFHsNBP+GeYdPpSYR1Cotd6uPtf+wORGD8K/IAWjr3b5DW500OZniAH+gk+9PE7gPFYheJgjVFapPhtt2F3ptJ+jtW
bdsyKDY4CLdh2WBXhoMBDueQXPKILzGPaAcv/lylEM7NKqfYEDHp8p6S88E+cxEIyBcQwygSjgODt4CzbHkV7411SZs1WFSHDs49wVBhU8wAF1qt1WJJ/LEM+4agJvfD
TPQNXu20s8mKx5d7hT2HaymgJyNAvCBfHkB0NmLnlx5gCnecd+6kun1o+BnpYnx+Y0MkFwtP/zh+P5KJZRMV4W8qXcYZILMlvVQE3/kHajmXMCDc25OiN1PjAaUxfcOb
VxBcZAVcNa1RS7CluMjjxEXz5sQJqBO9wBshd8nExEuwjdCGxT0NrIYAdhynzpfXU6dJdiWb2tYWmSuhni3ZmSmxymvKvkQHqPgGJ69+NRQJXVFa7Ppte+dUzFWL6CdC
nqXj3Q/wFrABYLG+ZeyiWnoKvmdbgtnX+hoZebQ45NGhPFBu74odqS/Da7QXSM+yH7qsns+3drobOr+zOqQIWy+JJLty4F+gvYtdv25FGjIMYaNhJf+YmFRl0wU/BmPW
5kOXmFgo+6pE2K1QRm4yAxnS/ll6939QW+4P5q4tSXZNAfYBaVa7LcAxttYaet/vSgEQuSBNhFMpCWNGJR8ChZjvqLsU2pnWmUMk7OfTFeSCduX+QcPi7tW1UD1yFSPE
zSEzcELRp+EqbzXJZuw5HNF+rhmdFSrwy4o/laEV+WBDZqTxJ3eXNBPaYtZA5k5YVOQG4KKWUs3uPzmlb977gIC9k7oGCsGY2n43lTnFQXX/1HQ2S7REcQOKDEBTsRry
gnbl/kHD4u7VtVA9chUjxP+z3xX6SOw4ewPcpv3/PVH2L++ZOnNfZUhD9SVqHqgZ4osM8cVwGLU/LJ7rhNRrSxov3Pc81fyEe61nDfnXLe7AFfExCs//7Qnm700GDjyK
vqHZtX0d6u9maEArfsss2hSERk0dXfq7oi3zCEtMTgKIB2W6U9kIgJvicv/N9ClYMD37H1E8cVUgUev8YpoK39v5AiHFH1vvyi0kUwhdOmMjPlTJc+aE7PSzruqztFxm
bWw6FwO4xaQXs418FVxyQ4l3YNcqp1dfw6l5rgQXh64U0tFJPseXygklEunBjD11o8gkSnokMnwQx8iGKh7X0bsirpaWCUna1KqxBnrw5ur/nmM18mnK2shnGsP5sGv/
dmMbHdMW/tRki5G3Hpk389ExUp6zZZCEY48wZfPIcT3JJIQXO6S3gyMBxSvJRLcRGbGvRNVp6y4KjprtATayLba+78ekv9QV8MftHHGjyi00NBM/cpEPrKcgq0k95ELZ
m+AgNlfnXEIJkn9FiX4ajLUW1NKJLB4LT5bDVGGzIJ+u9ysH4sn1wSjRHKQjQcUfQNZUdjXYvdo6L+xLRXYwWLxEsiUaRqpx8W5v3Ar+24AXwy1p30UCYENa8PYl1NH/
IeIg8YZdnTAxePyaHru/zf+Se8Ebv8Tnrw3IA4OHAGJPWGL/jz6iYjkjPlpeYKlQ5ROhfSXNFHm8+bHB7URdTUcuQWL8VUWKOqV9t0cIJdeqeTgZ+SVpiOsvCyapeI2m
yg1AEImUOwbQRw/ylC04NsrsV2J0jruYZwZNHmzYcq1WyCYaU4mJkJJ5tszcE+UkklY8lYGfULYg1KKbNyhT6fgn/78XqlwfPhr81VIcMdf7j0PBEMk2P8v9GizxMvkF
HRk95mzOalKNKksFARHB5SZEO0doZMb4EcS8Hr5kaivk8m8KRAgzTjImwHxeE756+BYkApL+aWVvAuh0ecmAdNmeIdzA0QgxI7QVzFtsN3B759sBdrFn2JYemxhxu6ae
F2TxROfq8uDH6w4kHDOr0KVPYxtrPkEBupNLTPhotKdHLkFi/FVFijqlfbdHCCXXtoe+nA/G9igeP6lrG+nA+wHe9CcQf4OMUuNVz4UDsMsYNxVo7QpgWEosKSjxAMW3
6gJkgjVMy0Ox4PTrI/Dne3nD1isIaO5zUkNHdWU3ApqUBfsTX2TDPEcvAUbZO7pyvdJdYdVeYxhVWQobbjKXMcNmc3UFc0W3JT0qrdPVXprZd61eBucPwWRqXTUd7D7V
njbPu7AKHsp5dIDJ7a28WriLl/r3/g64GVbWJ5mPmglsiO0bmZI6m+sOtpLeppw3pn7PSelYkK1URikSeIt3ZoHHQqJm1MI5AO83C9PRct3Wdj0vB9+gxE83j6+UP2C5
Gpp1t/8eE9oZgk5UhSN6nJPXhcaBpkDDlf1NEQjSp/gT8WA8nkIX2iF6pgpHIt3CCUJD3kCF58UqEvFR2tElL/l/4Ki9wzgsYXvFRtfdh2E76izWqSxCIHy3gEbUQnwq
NrdMQwYWxtBVgdzW9+lBITMn/hcDf66WOLqsuCe3L/QGnqf9a8oXQ8r0iBr33n6bCUJD3kCF58UqEvFR2tElL4iT2w7+87rs4P2aKbXii7Dgo+jSVYuPeOMywRCaMNPk
hUj5875ZK+q5ZefwBEt5hndQI/5vW3pAEDtJ7UoGPAOl7TmiTMa5bpauIWOP7hzmHWe+cimCI4LoAxuOP+txxs3OqvbosFkAM/spQ1QrRbJrM/PUkoi5pQ0cSURGoJ2M
q1fNZUwlhQc38s3KNghadkMPvIx1U3vqyqAPnTIeSFGWnTJr/9PfS2jsaIIAZ93VVfTzGeE6sjM6aEEWhcTrgwFeBog9tG9Hg70d094l4//bLYyPDHzB/v6raV2lwSZz
04whBKcIehW8/C0YNG+CGvc/zBj5IO8tpdIUiv8nrfFkIgfPBWZPyopI3O6XrcWQGMKTWYvfmikLz8ikusdHOvfWVPSHeCpGI/o50UtVnKn/PMD0yFXgRZX+M1hPqsKD
u5UHQhGqr7XYEu54Te7Ds2ezJFf8fp8fIRWqWHTpMDl91qZGWsr9bEr0GBAxLCV0QjLd4189Ii/uMMnufHl3oXyHPixWIgAWOGUBec/OeZjYHkhwdcaycef1mFfdPRGQ
T6Z/ZeQMOGgudhSLEaTWClPPSxBcfcxVu1XdxnPQeUrkFvyzwSQek46AGpIsETxp47Ue90Y+g/h0xgK0gLZL47D9nqFo5F6JyaVrxqGKp1NQsIRnbq+86r59p1VtwlNM
IGnzIRYbh259ovkXortZrM/j72x/jHGmyJpw65ySO9Ye8TAkIeHvsJg2vu/BwVsCN+P1axQwL3rBI34kaD5AxbN6czQeXN3nWsKwRMAA0DUzb97VBey5NfMuB01Aa8Ij
zL1Y7Lg2qDpBKRNH1WPir5wpggl+s4u5OVBgSooKSKDeCPLm6SreyCWEsFE3hty8Utm/o1JJwghf7H3y6zdh7RijKu28OnMmKgUiz935ZUQ/+lUI7lST3R9f1X/w0GTh
yu+0QeiBLalTkNhDQR7LcdjkBSZovlqRxLySWAl0mQv/74Eke8mUMOskWZXuNwJToF2WrEFlD72TLEf3H9XwrDFqWEbPB7a+O56BUi2+HiTfql9fgt3f8oNFGv7sTvy5
IGnzIRYbh259ovkXortZrJ+GQB4lCpCQUjKWrE5JJoYHUOxEX9PHYe7cWVAfM7k3UD0BwNMgiDFqZKzWrBEXyqM+9hqYUnwCwWJEAfhpoZ7Nzqr26LBZADP7KUNUK0Wy
uyoHZu0D2gDG7SnWnH15ZG9nPxYcIBZu+nGsqy4SQD8H+nbIOBkQX412T7seZ+vVb2WlEq8LTUICUTetZxteWoJXpGJrU1ZY+t6574RPaS1TJYSzXjGyWzdCHnGLSmhd
voK4rmWMxT/6ufjvKnYhTmBGftxdlxIHtuizMMA8vyQ7K/hSe9QxJdN541DxzdpcfIc+LFYiABY4ZQF5z855mECv9+r2sMqZS4tOxdLw8Gtk58NvRg5mXKM7i7uZVmc2
2YNLzKCKPjUtjfcfghY7c+rfSpepYV7pkiMqxiIm7gWeYWjzdzwhrNDFY1tx3p28HRaaM2JTqeTwd1UVA0G5YcSYE9KTQoJnkpNUEuMBl4FXSq2xzShHtfTptNGC6v+Z
WskOKl72CArpMXDRXdufB2NDUcVBDbTfs30+lz5hTzkIBU7KMDUTdb6pMSQGj3NxYi3sm/FYkLOL6+H9fUUow/ifYfiqLxgTAmEGvzI+Tvcq4dJ2xGlpdhPfaqaRpcgy
J+3yePOgtl8mSNUQDcZSih0PO8KM1PvuLY2mOQA86bw7CgLIXtLOmpia/h3v5OwFWAX0aSq8jdPnfYofg3WoHQx2kKBOqdgyqGKhGKOdf04snEnIy1FBc/kNNMIolrgK
5dWIQeFu4DCLJTVajfUwu2Iab48ajqcCuBtHoGQzK95YBfRpKryN0+d9ih+Ddagdr0QmjCn2/KtuskejV8wFH5dIu0ZRrXKeHcC5vx3/QQMvvMxHPQdqp3D+diNDD5K4
qOeewx9zENxLwyZfLra4rkAyJqKGuEC8c6kSafpyw5aZ/5OSRoYXCtamO85qqoPllcwqvgNSc0ZYb2cKPlmgLTfui/pEOnLC71Vuq/6KDdocBjPdSXu53UKCToQUlTvn
OwCdrHBEfn6mb5lS63TGoKIH56/mN+Of/D2XL9C2XPT6yabGGx+A05JuzxosX7c5m9gTYeeU0JPm/IMCBezRaen3vTEiQzwITFNGpMR5FDlI4/3x1nDr76x3CbB3Zoaf
5dWIQeFu4DCLJTVajfUwu9Cz+iwh2XuSDmDin8aJezDQKurmGyeU4mxUkwAjeai2FqL6ozc38Fa18fy2vxZM99m8yEouZIVFjt4/n9KWqkp+mGZK9qqCi/xokH6xDdf9
DT120NOwqB6RQN9fVAgBQkogazM7L0oI5486ec+sUNGLJ2V2PvCiEGEO+KqrUptQJ1WBlhNy/fCQSCTodMuK26L+8sBAYnDeYAF5dFVjshI/Dct3WYGhJ46Rc/CnNzPB
bNTyQhdZ2hWpO0d+bXeYDxxZ0c9jEHXy4ySPUSaCHYUufH9sXOILPNS2aUZZvnxSlbd9eWkKHkLUuzGOzBgOG0YyIQjtSoq4mJVlRzMkA4i671uC/C/xktzQ2NdYR8MM
zc6q9uiwWQAz+ylDVCtFspIhARshWwfeuMs9P5EIl4p+mGZK9qqCi/xokH6xDdf98/encPFI1MNklNwdwhac7ZNN33Oj2BdpzaKaV9WGQv18hz4sViIAFjhlAXnPznmY
/dbWsrWoV2TLHrlsVhCMBcSYE9KTQoJnkpNUEuMBl4Fv8a9hcwu4qBfQ/TlOtZ455ty2UEllo+2tqkYoPlHwnG1Jo8rsqYuvDLE2tXQhmcHLuQgaazSeA6MYSDSxwfZG
xJgT0pNCgmeSk1QS4wGXgTyc1hfKpU9moQV/he8h1bN0Vba8oRKwpMyiFUUvzAq7oDWdcHYAqL0XRLFzTIWLTBRPta0wQD9cVSNNLsY5XDPgpTylGJBiRjb2EjcXt0yU
FqL6ozc38Fa18fy2vxZM93N57Eco7Lsb02brVb6VdmWVt315aQoeQtS7MY7MGA4bgWnudsqruPBnEeERVHc5GsMuZRAY4OaJPrnk63zH+B/R37qdzHA/b9I3x6f/Xfm+
tNIBchKK1fPasa5E1YGuPXPzkoY4J2AwZxy4yEkdqpGBfhlLJwQB/JSp3lQfz/5dhukmwcTmZUhO8vsOXysAFW1Jo8rsqYuvDLE2tXQhmcEGJQwZWg+hBOGXCsXypPhh
UOFJwZAyKwEwZu7HtI6lfCLLwxMrtW9oDHpbiHkif2ZAOkgND7ZOU8xvSPrFjZu8lSXZ8lPw63vBEw3Zv4b/m/DH2PFr+ghQUtcfT+nHX1WpW7oydoEIzKy5bz5sXfa0
kJe0dRu9ydSsdAOeehmyjh0RBSMEMES7kzGbsSya3+GGf8XRnj2ytCIdSNkBW0pBt459Ul7tGICquGPrRU0aNTypfabJGpLdTg5hAbX1nsBhuKwncgUKvQUo8l0Mgow/
V63ceEQWzJ4zoyj/cFo80H6YZkr2qoKL/GiQfrEN1/1VRlCe5ihMZykm3bANPuaqYx1WpJG7WD/Ii6RtrJWMeM3OqvbosFkAM/spQ1QrRbIgBaTSbrXCWvAu9gVRV0am
b2c/FhwgFm76cayrLhJAP4sdUtEuSdZdPKvvwQ320MlvZaUSrwtNQgJRN61nG15aHFnRz2MQdfLjJI9RJoIdhXIJSXxDDedetdH4JMkjtsYtKa2m2zfMwXWoCkAXTqs9
Rgm8T5j4ftI3YK3axnR+U0jGwpX1xVupz3pPEAag3Qi671uC/C/xktzQ2NdYR8MMzc6q9uiwWQAz+ylDVCtFsrEqjaf1RCsC9gLisAyCc2/4n2H4qi8YEwJhBr8yPk73
X+FCdPtWVSUCwQ5APVzJ03gVRt0RGzFVQGKmeAE4aoIw7xWzt/i+oKWQ2eSI750vX2kIECVWqsfaSyL0s4ylwlDhScGQMisBMGbux7SOpXzQ5lfpdZziNvOhVjrj3Ma3
6Mlj+wf9dvkA6ML7EeiuI1LHolebDXbIldxnP5shBNVew/spISvhOyHjM9AeU+Mq4KU8pRiQYkY29hI3F7dMlLqIOBRwkE27a93xbVamnCGIxHUJM5ly5+qK+nd5Q8+q
UoVFcKVfDxQgIw11zv//hmNzPV4V+pUi3CzAZgzSZlc1vuMxrUMLytV+4t0QYxECRgm8T5j4ftI3YK3axnR+UyGp/NT2hKgPDpiDEQInaq6wv6XmLGaU/dbkr6ra9uJn
hwSytH5vFPefVmBb3qXAYgPBeBjTKeK5X7CstGnFvJPG6sb6W+ulySnSp/E0BIwtudGcbkpGp5Oa0gT4fOpStlDhScGQMisBMGbux7SOpXzQ5lfpdZziNvOhVjrj3Ma3
9xjUzK9GeWSiuRt6gSZmlXEGdxDyxL4mAqzOEoYAcs2HQghReofM7Kouy9ygN52DWAX0aSq8jdPnfYofg3WoHSOoV01L7+igawnbk4+zTYYOTJOdOE9YYzho504Cm7hM
OQn+z27saTsf5/vBGJysxu3XsZtTCVHJ0AWd7HJzLsVV3NjcSLDCln1Kil32RD+ksNrRM7pVU+Emssz3d1SflEld+teYumRIBPsElUMeqzSoD3kUooogUi6zTOi/6Cb2
XFf3lnOlleeYi4vKZiy6K1gF9GkqvI3T532KH4N1qB3iyN43iNeFvHBlmcUGHUm+e5vuWQDgXqv3Xe9jHZ33bmuOQEBPgr0W7RC39cz56aKc6qdgiyRCL2kN8w0PhI0a
WAX0aSq8jdPnfYofg3WoHd0q9JGdi89VfxM6JuX46xzK386dixahGMyFteGR6nl15MTHwCPNcns/aMRXjDbE3nLBBuVDGY3aDNirmgZIhF1HbE8R0jHvFGkRAPbPyPGB
7OA1z/RpJeLZXrOQM9KavTXFZoM7604wW7FO18ZpACjCeGlVO/DCgmv9+0YTEOITW3ayKvr+k050Z3ZVc/dYb0oTqm44i77AEPZCg1SPKk/KhutP56KtseqsBQIPMSVz
PlmmflFSRLdZFMj6Xp+XoB5PJL9qP+vQ0Ql2tyFYPuIVzfG8053+uTz8HSm5n0GLE3HIbgahy1s8Uq+Hv4XiCr2Phv7ZbKtCltOima4yArr85NHpnDmBuD9NevsJTAAM
UnRZ62PPSDraPLbvRg0s7ZDdT2rcUC5+gEQ/BhhH+/U9RvImJnl2SigCuaqldfj6mSIblwn1Qo+Ow4rtozjvs8J4aVU78MKCa/37RhMQ4hNbdrIq+v6TTnRndlVz91hv
hsUGL96elLg7ZkVlzJMG7lEN0XFVS7qPH/APwydBTrEcJw3uxYp56JqUmgKikT4tT2o1pp43hR66dx0kmZZbwaAVOgnnGAPZpVR+7Dxc6FNX4dMpzvePw1iW/Hg1ibFy
w8pC2SqXiQ98WH/Q6n+MNbMV9cGuDeM7/d+QAJ9y6+Nk/UnI/mUEBVBt5SL1BStI2BvOt9oWbvVKGteVSSjcv3xG3c6G5nHpr2kZe0DCO5Dl9nfpk2x45uphsZH+FecA
adQHe9rZNvBVfeNlmdsWnvvjB7CjiI+nkj+VhCBoMReXW3Evodw47Fs88IbftbC/7PM6cbzV9ZpRfb72bmTG90YbYoIfGMlocnCaHag5cC3C2UjKH6yKRgMTL/U0QH+T
knVfFikngIHMkgsguEwex/BhdTllhwCUREzoGIQqWf9DWL6V2aTEX8L0YIhZC/K8QtkmfEUtH7Tn7bAuZn2X++zgNc/0aSXi2V6zkDPSmr1iKEX/waoKjY89J4gSbwcK
Cgy0NKkAjaL1LnsSPycgeVt2sir6/pNOdGd2VXP3WG+U/AebkOF3RV9OvtAQeliDx34QhqnWLz+iY8uqe1LCw1fh0ynO94/DWJb8eDWJsXJ+aPJiyn02M11DqOYuJxkN
Lby2F+TmGpQR58qPD/+qlzIoYZK+3JYDplrDcAkabD29tY0ljp5MfhyoNEpJna5AA94Zyqf9REzG3RXdUDRDRxiD6SSHnGWdYQBL69oCqxu9tY0ljp5MfhyoNEpJna5A
A94Zyqf9REzG3RXdUDRDR/F55KdoxXLkxdncoiPJlKPr7YGHIrBw79ZVXMMfc9jP6bxDDJTWZweftMZenkFzbxyVCOaw2bgjbzgxUzUIqfLj/bkc1BJx03iblosxIkFM
I1oyjJK2CDhVNBaEqfAXI0T+BI8RndVqmM5iLOUO/VKnTRtrSO38MSIrkrYR7rEvifaBY8Eu2if5/OStwVXCgCR7bQ0pNUVUE6dyqUSD9j0epRzzNXw7fnFtOimhdQxA
R2xPEdIx7xRpEQD2z8jxgR6cXQr6b1V24SQngTS4csnkBuV7VwjVY6ovRO3eB7ZekyjNbvtloOMTsWlhkUC+Sh6cXQr6b1V24SQngTS4csm0wWfOC7LMoJSkw37A51fZ
Cgy0NKkAjaL1LnsSPycgeWvb4VrASi9PLx86+c+9qEmHpAoWrnLxqgG8RmKW6PGfc8UHxHczZzqBg4feOXkHi4gsTWes4dfsZjrqVIdkjINh8qeoCvSoPu0hYu+c4nl9
DaoT8A/UVctujU264+XwRRpMfELE67dhgNE9qMs23vfvwcdXfPpo5KZWn4GjFN0mSEA4YtIUX7zQF6//FAyfF8LRmYRNn2qhGStGQ7nT0RWoD36li7kBGH+luCaitgy7
ifaBY8Eu2if5/OStwVXCgGfnJcDMYunsPdXeMUqtu+1UaGmtH5jOqD7n2QOtf1FI0m01UOOjYLG3z1w7I/GsA2fnJcDMYunsPdXeMUqtu+1XrQNMK5QwSnyaBIs9bqVc
zA3Lr/3Q4LLy7mjIFCwDFQzswQRgkID462YeVL9plHGrRU10XbAqFT2AH2j1tdBxzA3Lr/3Q4LLy7mjIFCwDFQzswQRgkID462YeVL9plHGCrbG4jwqrLHn6f8pOCjr0
ORmyfQQVIsDj80WVZb3fwQcRT3H674YbW0oCA09TB1XsBgGBZlO/TDzymf7c+JxleguZZBabphTvYMUapSttMllTb1jCz3INO5We2dJ5b3+9j4b+2WyrQpbTopmuMgK6
NV47cAtxuVZoE86JC/Yh96vcPTWWEGkZ6nviJy9wJpTjcJaGqYdvjlOod9sm1NoIjWtTl7bl3NI8Lkv4CgXM9+j3fQbjy0X0CWRe/Bjcrretlj5d1KQfiVjqiZJJY1NX
mliyNTbqo1vWB5E3a44CN+6grcv57j6WKkylgZSHIL/CeGlVO/DCgmv9+0YTEOITa9vhWsBKL08vHzr5z72oScR/44dZm0SWwtJOqbqewSJgg7vcrtG96no2iycQj96B
T2d+SChpd49N9Npuzo3d9CLT9m2c8IQM4H2ZXrlLbIQLIfur7jh8WkxzquW8JRALuFF+e6TVrsoC82ybZql/8EH3xnBHs+Anu+hgJZ3uC1egU3uAd5P5mx4yFH6qOu0i
JY4rMzP3eTbp2cvdFKsfcasrkM2tE/PoUNncIMJy0eR/4EYoPUyDK8jVJtxEk3EWekwXK3JLXctUs76x/LKJ2qGNuihNM98latsGeoB2ZkwGt6oyLQwhyKwEOCg6SnMR
/MyrXKvn/sN4bGr25IR3TGOLKN/NVM9esVtn30j64slFTtzj4ByygKnyQoSrGrIy5/jxF6eA+GcZ8wZc5uJi8oRluufNXCcvXBa6e+442cd3joYKtcc7x4wCUefzRzoc
0vZ/C5D4uxV8hGR06yAxc7joFy2qShaGoxPGImWTJY5MMqO1m0a4ugAp0OuO1l6OnzCjI8O0AqAYsJaaCTXpDqBTe4B3k/mbHjIUfqo67SJxffoRhWsh83/AOfjTqRbp
ApA6ufpI8X6/LKIymL2NmaFu3gyTYk4hcryXuKtshg5yBy6pfPxUoXEONUlR82N2RPSVlqBUKpiz/b3JoD4gIBHQo4UKRp+0DH573OLeJa1sOb14VGDT1yeFC2Vhxftz
Ms6Yp83sbEijSPVFltsRMEVO3OPgHLKAqfJChKsasjKWo8tcFWt5SD/7ZDqDO2RH10JwP06dEfOFAx5dqgo61JTQt7OWX/w9bQN7ubvgcLfS9n8LkPi7FXyEZHTrIDFz
AhB7UbTWe27yYQQH7EHcjbhRfnuk1a7KAvNsm2apf/ANtRGuwj6Z6Fo/rOyHcVqcoFN7gHeT+ZseMhR+qjrtIh+ZvrJzt4In3O6CuYs5KY8SN0i7V/sQLVUcKVyaLpFU
q62Mr6lg8nnIULcdD2QwCXIHLql8/FShcQ41SVHzY3ZE9JWWoFQqmLP9vcmgPiAgoQEGP4pjJ/q/Skw7jsGKyjs767iMvfBSXG63huhS/MRUxpQyd0HAX6TAySxe+F5G
RU7c4+AcsoCp8kKEqxqyMt/T13w2knQq41DaImLwW3ZRdLU+MzJ+N5nbqR1zCNdpoB1H7eess8hzaBA0sl1vHNL2fwuQ+LsVfIRkdOsgMXOZYJulv/ivO5Mecm4CJf7+
GYwcN6DmUuh32QcbDRwuyZlgm6W/+K87kx5ybgIl/v7px1X7c42EOenspv0DO9xCvF60JFPiJ1CzyMDebSj+moSR9VnxyDfdFk3n8BkNSelMv0CBUdssLJrdUdYWu+AI
cgcuqXz8VKFxDjVJUfNjdkT0lZagVCqYs/29yaA+ICCMnrLPeoffoqQfSlW4rAPyBVgSdo2/fUPtFBGp9Hn3+prScC2zplgjK6h+57ZKauRuE8JomAdCaF3g9Zf84UgZ
7faTFUbBaPxeiIyrHYpsAOphpReRwQzrtkbKXZeeUOszzoDMOLfCdOEXTcrvuqJdql1NB7U/njFU5faCQY2X1xEMPkgtFdUYaBmyt+yGjhEZjBw3oOZS6HfZBxsNHC7J
JsfOjaOJFCdI32/TV7TxM7wqPJy7XgIJNPNeKFZpNgqotzJ8kdoaEKOUbaa+Bbj/x5u0YqVe4kSPsanIbJ20e5PHTDhN0lPFYtfPd+ziSt9pqfkNMYArugGWNCjb4K0h
BgFkoZbbTLQ27IEut7gPkfeCgDbrD6K1SWXtPrNbLSpX4dMpzvePw1iW/Hg1ibFyb897HZAWYDNpUZ4Zvxa+724TwmiYB0JoXeD1l/zhSBmnsYm6pFo/DxYVzEebSuqQ
AiTFyEQFu9DAxiJzQEwaZbFSkEQchg0CCKwa0FlvnOrS9n8LkPi7FXyEZHTrIDFzQjOzrklLYrT6MfUQ4f/U4xmMHDeg5lLod9kHGw0cLsmLNWm75OEBOysa8F+kZnxi
/BRJMnoFFLKiT4GGu59IKFKnWpVZLdoyP78eNEGSL4we3ql1ORnVqaZ0LWctn+JPh9OA3FLJNvfotF437Fr7eyBpl7nzuKvNNskG+6HIXEIGAWShlttMtDbsgS63uA+R
DpCOo+PHHOkhi2tXjkq++1fh0ynO94/DWJb8eDWJsXIIo9sMLPpF7ZCCeqWOet9NbhPCaJgHQmhd4PWX/OFIGUYe2bWug01e03nwprrFus3qYaUXkcEM67ZGyl2XnlDr
/0revoJPQJyh8ZJLdVI57apdTQe1P54xVOX2gkGNl9cDJp1PRhagjMEBbd8tB2uMGYwcN6DmUuh32QcbDRwuyRwbeo5kEFaFew60/nvvzgZue+SZBkZNm8m4v98f1nZC
nXoEItr2e0XJeJoNmBJemk24iikmN4yNEWPFN8nVE207v/zSiW+mtX38sbpZCq8mvz93D/wsdQNPDRW6vxXZ6gYBZKGW20y0NuyBLre4D5HRnOeM7tafumdu4nEP9iec
V+HTKc73j8NYlvx4NYmxcgnU8esO06q6216U6QanP6VuE8JomAdCaF3g9Zf84UgZRR/sH6t8JKEmzYodP60c5uphpReRwQzrtkbKXZeeUOvHkDgsSXne1NgGX0XFT+oL
eIJSTMxgJn4+DLS+j60TU2/DuiQkAxvFIbEiLlh/m7YZjBw3oOZS6HfZBxsNHC7JiYcr96Wr4B8rQka1I8nCVLwqPJy7XgIJNPNeKFZpNgqow+tA4MX+NBAlq0F4VCA+
gyy1q4Tv05d7xBLEPVyQX7UShdSWzu9bQyokay76SmWD1rGsUMNU4oi9/CgEJ+DvBgFkoZbbTLQ27IEut7gPkUGiXPQdhslrE7r/8fE1WhDx4U0oUl6i6YSNIlchnsCK
yogm0Sa9h4GMq195YwJtiEVO3OPgHLKAqfJChKsasjJo4J+ge0M5FEb+katuyyxA6mGlF5HBDOu2Rspdl55Q62jgn6B7QzkURv6Rq27LLECqXU0HtT+eMVTl9oJBjZfX
wS6UQp+3TPKF42QeFPcvmp+l2H0vFo/iQ2KucjogItTdbSbN+qEmf4gecmKn6DZ0oFN7gHeT+ZseMhR+qjrtIk/ELOVTbrzyz+4jUg/hbsxgq1WQ1al/4sEkvWSq9JaG
FktDBCYb4tM1WJjrXeCZ83IHLql8/FShcQ41SVHzY3bMlrA6kAKGmalSZre6myAH94BUMbz8OQNkgU4U9TpW/zR+nPAiirPvW+brJGnN0CZUxpQyd0HAX6TAySxe+F5G
RU7c4+AcsoCp8kKEqxqyMnI0KrbmKFCVY48Fs2XrJCXTf+NplqIwiyN7cV/azu2yLmKRiI2lIu7X97POMWrj69L2fwuQ+LsVfIRkdOsgMXMVCC53l7RTvodGpy0E48nD
OChwhrvOT1+LtITHLffs5YiTzaeBQzdz2bF8pd5cNDKgU3uAd5P5mx4yFH6qOu0ihTaSecSzk4KTTipR13FgHySSCio3JmTYuwiVbOYm/cHJ8PgCLzYC/VqdgpdS9Wsv
QiH+6sC7fVPv/ZRtl9Kr4zbr1KgsfVtk4fzCsz2rmnkq0BUiesPcoBrUTtR6Ks8qpuXsS8y5MoVI0/oDlBXdiQ5Os2BW18ejZdkopZ8kbUBYB7BzPZAKE3euKokFEjHo
uGFo8WqpN/a6gxkKh7p6/dp8KaxIxCfwRJJPZaJ4EinTIZGc9kTWzrYMDyDvnYgc80s1u2OqHYTm0Fd/2Mp/6N4dUnit9vxzk7l/HYQFUOkSOZ3Kli6K/DQZMQeKYcoA
f1YGlLULHLsY6rHP4SzBB6GOGRbTFlHiOvUQpjJMgs0/3HRTH4ZGRADEKVwAPIR0WrIFbJI+yDQ9BMRwNxmvM37dAyFF8Y/sLLa3xBIpOrkyzpinzexsSKNI9UWW2xEw
9rswH5Rl3UkeJz+f63rT7/BjdbRdG+PATe35cQtL6h4U4Cct5o0X9iaR+3u1mRYA3+g/XMibzkckKX2QO8txWcqIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mF
sb/kWnu4Yztq4q/g9gtMabhhaPFqqTf2uoMZCoe6ev0uT3tRB8ZsijyfwZjo8FOu0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+jYQGClf80rL6Up9Q2D6Shv
HGbWyG7K7D15UO6nQw9l9R5ma1MW3T/RqwHknG16gBeeQ8QsxJAEjcphVGeA8TFGP9x0Ux+GRkQAxClcADyEdOn+4eTokvQ9tjW44DfiXFpTPBTcMRwSlYjDZGMbALTi
VMaUMndBwF+kwMksXvheRva7MB+UZd1JHic/n+t60+83a8UZRQ/UlthJIsdBxcUeW54Osm2f5fxnZBcx801jQ6duDZ5lsPpCAJElxmMHedzKiCbRJr2HgYyrX3ljAm2I
bcx9A3euJafUPZh7l1vZhZtEAJdlCaKk2uhuCMLaOsu4YWjxaqk39rqDGQqHunr9pX4eqdrWKSEgDnR2v4/rBtMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o
tmdT5/ac/Qgg6QMUmBN90zSyo0W8/Z4+LI43vsp7lYa8InNUSLt9BTWEmpjTEYlHnkPELMSQBI3KYVRngPExRj/cdFMfhkZEAMQpXAA8hHT/5kZMaZisfWehxUOgVy+d
l1TgTWvMurZ3y1ihSz5NdG49yqOPgox/MoPbrhsZmZ32uzAflGXdSR4nP5/retPv3frN2nN6gvofWonKf6Mx/BTgJy3mjRf2JpH7e7WZFgBqqx6vnMqFlrrXP7q7NnwN
yogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YUfHgL87WsOilq8SczXnTHViB87cF+ADfzXvjg3uLstvd33cmDSk9SKNleh+t8ICqHTIZGc9kTWzrYMDyDvnYgc
80s1u2OqHYTm0Fd/2Mp/6DAjKrP79fbP6Ik2gMlU49sSOZ3Kli6K/DQZMQeKYcoAh5raucxvQrsv9VXSpUd9X6GOGRbTFlHiOvUQpjJMgs05NRCjTWDposRMWfMGo2Il
+Zg81Nnl7bouzkaYMGoV6PbqZ4rXOD9atMwbmK4n4HFUxpQyd0HAX6TAySxe+F5G9rswH5Rl3UkeJz+f63rT723HqbU35ondo3B1FBZt3isU4Cct5o0X9iaR+3u1mRYA
IxqDFtXtG67KZsJkTuFB78qIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mFp41byGH2irnPTSLHGq3BqIgfO3BfgA381744N7i7Lb1UnYDYG99HjGn10FyEDSBc
0yGRnPZE1s62DA8g752IHPNLNbtjqh2E5tBXf9jKf+iOXenBtQMYYzDihO2Ri12TEjmdypYuivw0GTEHimHKAAd3wz85WIFf4ywLsBTSLyWhjhkW0xZR4jr1EKYyTILN
2C9MjKSoYUkfyiJpguDYMR3XOwv9AxDxLTW8bQKQsfF3TGXmmjBL86lV7xae30Wgyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60++R/cBM6KKvn1LEMN8aVxaY
qEr6N5BasAzSpKvI3L49bTHJWlrHyAA+5mguLKecKT4mEuSCm65WyTiOtqiKs0/bEkaolafW3+oauiKYwUAYVpqZUQOsO9peVdKN+KmU5nCqh4scgrRMCxmN2SgkPFzT
6iSDJDYdv12K6Gc0O76GlZaQ5ok1rD2jnlRJy8CxKO6SNw09cGng8UC0zuarcnzV9v8YkPZPC/wAc+pzSxkrthI5ncqWLor8NBkxB4phygArrd+7B7GBogm4HO8GIJgk
oY4ZFtMWUeI69RCmMkyCzfu/eVKWNcYmBrgRFUSyqi5P3yzaNu4G5509tai5SFAxX5DQjlxMvE6RupzNd6nYbcqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
nh3JQaHWKOEEZzc2XBAzg4T9KFMV4KE25XM/6/SaGOY+07djT8F1/avXwdvrJeYwUQtKb+fYpkoggaoOn6jJ0xJGqJWn1t/qGroimMFAGFYMk4KvCxNcAe8BQun27qaJ
T79LxMsjvgwBClgF6F2BonKPe+w6DKZ3YivWt7JQZz4nHskfB9QusOl2qjoY4Mx2kjcNPXBp4PFAtM7mq3J81a3QjooRma47KJl4X4OksTASOZ3Kli6K/DQZMQeKYcoA
JxXwIxNL/zvFOHmjMbuBznRy14IKvto20rLBjhPpzHn7v3lSljXGJga4ERVEsqouneipdb94X3kvbqDkHXtATMLRmYRNn2qhGStGQ7nT0RWtywArBa6dMsMhQctS6nCg
QMmqsJAIM6uAKSZME0akDBZ063V55GjuFHP/3180aRqE/ShTFeChNuVzP+v0mhjmTYKGrGS8E8BoU4aJw7+f1ldq8YsnoNZVKDu9hZNFIYESRqiVp9bf6hq6IpjBQBhW
hMtqEeg1I4v/F1CuZBgE+k+/S8TLI74MAQpYBehdgaKs/YBWiDioat9AF7XVBd2c2BndPvqE+Zj64oLGTB6I/ZI3DT1waeDxQLTO5qtyfNWKYSE2EUySIcMutRJpYIPH
EjmdypYuivw0GTEHimHKAJPAJQ3dkvW044/4qwkbguihjhkW0xZR4jr1EKYyTILN+795UpY1xiYGuBEVRLKqLgv6HNGEMT3iXeTD0c3xhZXC0ZmETZ9qoRkrRkO509EV
2VLVXSmDXq+0XXtVuFPuxkDJqrCQCDOrgCkmTBNGpAxnbtzmIBRXaT9bbQmSGyZEhP0oUxXgoTblcz/r9JoY5vJbMrv+fkVx3QQGlNTCYiEdiq6lKX8PmIh8vQzvhFQx
EkaolafW3+oauiKYwUAYVuJoCRHHCwjBxRQKeqo6IEJPv0vEyyO+DAEKWAXoXYGiQoN0ID83OCkb/qzHY0siIwApOmyYw03MoNG/8da6LG+SNw09cGng8UC0zuarcnzV
npVgBnfGaYE+R0bHnOQTcRI5ncqWLor8NBkxB4phygAPFsMfG8WlfO5ZfNu4sjfxoY4ZFtMWUeI69RCmMkyCzVucZZBHqYs7xAAnIN0w4a4d1zsL/QMQ8S01vG0CkLHx
hgAU4zZAnWmu5x0AYua158qIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv4lmFxGSh4hYMP3zjhSIqOYT9KFMV4KE25XM/6/SaGOYFwOokQh6J94m4oyjOYoXo
LnfpZMUMik0jsG/ygpO4HRJGqJWn1t/qGroimMFAGFZ/ehjp7BOjJiOHJliXdwJgT79LxMsjvgwBClgF6F2Bovh4d2iMMu3PlLWPzrHch2vBB/NfB0P+4TGXuKFbXtsq
kjcNPXBp4PFAtM7mq3J81RjeYSm2VM34dabATX+7JjESOZ3Kli6K/DQZMQeKYcoAWWT89wHFjWq7ekXeFpx6XqGOGRbTFlHiOvUQpjJMgs1eZBcin0oHXQ0fk5THS1Eh
FyertMzh+i6zoHp1hQdZCph1vWri5PXWW98ih6FtOzPKiCbRJr2HgYyrX3ljAm2I9rswH5Rl3UkeJz+f63rT76yPASmKalKJGkKRL+iUp/WE/ShTFeChNuVzP+v0mhjm
p+M6QBlwV0i84SyRtrdil7FSkEQchg0CCKwa0FlvnOoSRqiVp9bf6hq6IpjBQBhWjhBUmbNndoysNgpFTCTRQwYX5T2mEvQXkY5atWu8OCtzRdFWyTjU+n7mYfXaSZ3I
0yGRnPZE1s62DA8g752IHLnP5Pjl4sHgFuRC5wOFZuC3/b97tWwj+3ptV2A3DYtIXp5O+UfEMNEj/VFfZZpTHptDYAQigVsFfc6EpXG8sQ2eQ8QsxJAEjcphVGeA8TFG
RvNLUWgVRSDyLaqmkMOhGCaN9KqRKMAV+2HiwOPLtP1Yu0WX7WiEM8XSifi037E/yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+9telntkUjeb0MHJS6Uu/y6
QNuG1YF0DMQaoPi6gbKncjDNFD8gQC7qU++CVTMinizKiCbRJr2HgYyrX3ljAm2INR6toPpwucioa8Rr7WlO9DV02NtsHna+KpKaSs0i+/lA0d2DyGre9tvA3w68mW96
wJM4cwbV4A1gwzHbEqpRPBfDLWnfRQJgQ1rw9iXU0f+5BhKUstv5pjq4abBMW1/5l8aSLhUvhPE0T8vt0qrTD4A80proGFPQKt43RigM7grfMLqfRsVnV02iumKMqYKe
/Wh3OcEbZ1I4xQ+SzRV+RWldM3A8NENLO5iLQk3LAFVERkearOIYBd7U4KbAFklPzAFB8irA99dnU34r0QVpsbiqaRIDuuEKVcdSm224n+mZ2KZStSp1FV4bvJbSasjz
19/omKBRBEVt3ISD/+eN9uSRHZ+Hu2wUSu5F3uyuI4a1rM8D5tvf7watinz4jQFysCPBEkzfnkEUk1D023h1SoR+qSld+IIbqqnJyrU6tuIMEO691JIQLNtlUmUNWuk3
LBDE1F8aUiA0A1sJRJ/2ZlY6P5ANkRDrG6eNWtoVYXsbt8fUjU3tL03ExQTEdZtjqSQ3WEwtO+R1In/Ng2CR5Hb58Gif2uI0HXhyaYYRPIxQJgZcAnRSQG51/wte5N0L
S8xn/NlYimpPbSj0DP1dk4kK3ICywWSjKCEZgBY/qLa4qmkSA7rhClXHUpttuJ/pCktAz54q6+LbPBgeSdcEISbQXkn3wfIMlwKoYJuqo6dczEZvbSXWzm5shw281dOq
sKUlBo5sx1CAEasgv/DI63eGXjwSOcBUPWePG1NxFZ8m0F5J98HyDJcCqGCbqqOnHLeDk6/GCYhZxJmOCcmt7CM+VMlz5oTs9LOu6rO0XGa+AuVxPzPFnnYVHPpTg6wa
c0gi5IZdJqAsjzuYrOAUyRcp3jZLlQ1MJ1N3uX/RZcc1H6nOMZygF2+0Q2k4Jr+BV+HTKc73j8NYlvx4NYmxcjF0LACSJ3RpcmYKWuccjdSnhYytBVDjlmPef0I4m0dr
sS+mdn3hvPhX8k1EZ9Wmrf7Q8Vix6WX95uC7VWQJW4r5i3ozr+3XlcGkGoYSfaSNuRTnfisBS3XdP+g2JfLX2SUD+pS00UZRNBs26HnTLRA7aRiHyyAhBTD0bKMRoFJ2
ht5PbeBrhCFC1raSRE8TavnDbd5FoUmKrSXegidl01A1OWIIES5dTOECIF57l+fS178ZZQzuOkxWHBhTDWJ7HvG2sHq3qLAcxj3z9H69b4sRt3F9MrLiZrH5ZSsud7qL
L9oP1mYZ2jKURz7eAc6d+sK4fL/Er1/LPbXfHA5ecxnOKWl1u2/+dfQxJGzZkqO1HD7XwJRFP+IGc/XqZaAqChwnDe7FinnompSaAqKRPi0oFuLsQjNvffL0Bbtl23uX
dLU3k20GPfLG7Nkxe997PvK6jv5dFoi9GsNUKlLgbwhR7ZbTiCa3K3oPOSdi1hitNTliCBEuXUzhAiBee5fn0ssvzLouaWWfpvHILxrn0aYHuNIFTxEjpdqfmnsK5Izm
Iz5UyXPmhOz0s67qs7RcZmYmaB8n8BXv7YmVGV3Q3ojaw8o283qh5mfmEFqn5YfR3kVvo0QQo3hkHbha57RjeTDvvncav5NpUrCN+X7OBOIyKGGSvtyWA6Zaw3AJGmw9
sJyciR5BVQsqt42nTaal0pvIM0kFvw18N1kqcM6pbzq0OWdXekZ6+fWyLSJwCb1Ijt/cRcVsuk5J6p8WtozGLzpXyDxnySt5m229jTfXceOpK25lUpHGoddN/4XDXpTT
cbRStoYdEDWI2FYrIwJxLiM+VMlz5oTs9LOu6rO0XGakUnYGq4z5fJajPM5wxjC7hSggl8U9r3Q0UhRhjuSLiyM+VMlz5oTs9LOu6rO0XGaHtOjut1X9jJIlRJYugJgR
DOzBBGCQgPjrZh5Uv2mUcceEVokrhcx78HMid99kmgNJzJ6OtMWzDA6Xbj3djZHUtDlnV3pGevn1si0icAm9SAJYvdeXKIUrZ5d8twY3p+eMXUKaUQUG9XqCNvMK6Ccg
2QOppdttQjkEXVecVQJNJcJZOS8+nHDBEdGvk1e2C8XdWaSxAQrFiuiBmM3V7eGtJg2eZbqZZNg9AEeZZZ9cWsd1Ke45XDt9DGQkpetaiA7NVsFqNlty5S9rtCe67AJM
gz1Yld6Ng0NJ9FsM+gCmV8LRmYRNn2qhGStGQ7nT0RX6Bt70UYre5Ht2XkYD6audiWnXR0rGwqwX0arWVT7TGoMxFJLNZGyh57twpyB0yGFhFlHhlpF0juYsuDnPQpEe
3VmksQEKxYrogZjN1e3hrSm8Wy+y6kylFS2KDnI6xdMmoVYdGj2S3CVCZeAYqrdjIz5UyXPmhOz0s67qs7RcZplIGjCwO5V/FAxiPVVtIuMHEU9x+u+GG1tKAgNPUwdV
6941ZPFeylRW1DLda2JtN3ZAjtKr5FGfYDwh2yDNM6HC0ZmETZ9qoRkrRkO509EVi19g4z8bpOJu4H+RAgxixAvkuPoaMaqO+OdFU11rZ9a0OWdXekZ6+fWyLSJwCb1I
+R0IQRWqCYMww14kDXq7so80qrdX5VNNww6BDhxRaHGDMRSSzWRsoee7cKcgdMhhSFdl9FxCXnUxXjnnQxUfuhA0cRYQWHYQDQ3afcnMEhTdTodJYiTV6khcqIlcQq38
b7CRvz8+OKyhrKgRxPxOopTeZlc4ZkOWjv6US4+mJnx7fINgXTidLAjb+p+Zcu9m+v86IvPDBY+JEqxjWLs/FyXK0JK77nMoaEhpNpqE0FLbXbe5iYcraZzxjoCBwCyc
JM9na6twyOFbg41+L6vGwQRWYC3SxE6keSHezpglNLwf0gn4j9YetcG4jRrn9OCQVUVM8YorsMsM8rnfYwdhFdtML4SdHK529a+tCqokeEzEmBPSk0KCZ5KTVBLjAZeB
b0Rq6aBYnlKrpV0NOmLqEFnPUo7X70ODr4/1ZvU4mS3dKzQBErxYtdnAlT815O7bgEdaVG2oxnQ/fXlfSoGAgi5ikYiNpSLu1/ezzjFq4+tHKLmXaKvDVYiKuhy6u58G
+NyQKvxl1tpuRJRYhHLUUnnXfZhyNmNwiPmeZrs1bzI9SUvcULNVUmzeLxdtR2+NcohLipBsUL1t9gqJSGPO3TVgFwCgjHl7azLRiJpYD/mez9l7f83N4+GT82oLF3fI
1nY9LwffoMRPN4+vlD9guQWhApW+Fn2SszipHwjJoa55Ms0xsgooJJw6Ofj/UaB77cjcMqETPsC2d2PZiP0L5vg+xcpzcoORuJfLvBacAVIAivN9GllpjMzVdMrL5UzV
OWhWRavz53D0a7HZ+7oa2JYNGdfSWOIdKBJoJMwnN62Ku+t8sbYADGua3ezHvns96FJJzG66DVihUAr75P147fhrbHqZ/7HQjA9cN7VYwY54qVP4lM7CmalgcqIFM/7V
b9mVDeIlDzMdloUlyMc/q8vRKBMB7zvimCDssLk1sKwDCZrPdx1Oojg28ePRr9Hk1D7w3faJc63MY94iyxTRSdd+oxi8u+dzyk5VdeC8U5xkjb7owkbC60XvVJHOWzyU
fcm2hG+IOPXPFN/6VeGMmSft8njzoLZfJkjVEA3GUoodDzvCjNT77i2NpjkAPOm8Zm1d3MC3JOjUnf8H5vX+seu9iSp6hfStMsJxhHyV3tWQl7R1G73J1Kx0A556GbKO
T0oX2oSDfsmBg3GoU0Zq08oi8JXzLdmIr5+bIa9fc9PoxLK6MGnMhqf+v5PRiZ3zZEkljiuTsidH93CjhXspEFgF9GkqvI3T532KH4N1qB0SJHaANvR3/LgKNPs9OH+K
j54Ie9I6A2Eu1jlRp2uJsGNGIZ5FkzGoFcF3+igPZPLAHNOhlNYY/XL8cS9HF1SKM5Qr3qtLzEHjxmPJFnLZ/+xwIMQjFqApkD8SotWI7sHSgz5L/+96iNCA/Lyga13v
6MSyujBpzIan/r+T0Ymd8ypyDAfSnH2R1flpgIjDhkFYBfRpKryN0+d9ih+DdagdDHaQoE6p2DKoYqEYo51/Tooyoo4PPXvU0drwD3GDyKoH39EmOMVMnxKb/oAbdJxx
62sdUJBGmnwIAri7z3dXY8u6bpf0koypEhaaTKQKyZzHszVtAa97e1+EGcEf+MyXogfnr+Y345/8PZcv0LZc9EoBELkgTYRTKQljRiUfAoXuWMg+pnd4mpXUPbDf5Wbi
ZOfDb0YOZlyjO4u7mVZnNiNAfE8s1V0GiHixYgZ+wB+YiSZH8j6XUrFtLQy+6fJ4HQ87wozU++4tjaY5ADzpvE8U3CIBr2J6hNNClY2+b2YUHk78twSEGokH18AxreYY
bmm2KJRatMioOVi+uuW9zDzASfA9ha0yrDQvhqqd9m2wv6XmLGaU/dbkr6ra9uJnNTehDOFcnp4ec1all1443AbZhRxQk/b115uvDVp8fYvphJFZ6P5d8j7sxvrfevzW
MiMvU5T8ts7YHaviRNyHV7YEu5VV6RvRfKX0i2y39rtfEvePVOTK9912Q07u4PWdMO8Vs7f4vqClkNnkiO+dL0cuQWL8VUWKOqV9t0cIJdc7TEyKidjGnZhQZzkfkOdX
gFKh0E2u4dtRh+pZ+S3e3vsuz5XQBj/VJuzTxOSIlhYXbddjwSmIwa7XUnLpp/mbUOFJwZAyKwEwZu7HtI6lfBxOrdXUxq0mJ4K+s7B72YsYuay7vfJI6O3a4nZueITb
2RSRGFSm7XHFhiZdlmAk7aMjqWLndd2NuyBPaQf3NUTItVlA3/sRQe+PaLvyCQJzXO7hHnk/duC2aVOtdfWehogbC5KaMnWEtXqSp2Y4X05Q4UnBkDIrATBm7se0jqV8
GJCKhVWPqWAsY4KpVwW9qEINjqSk8+jzkcHX3yn5PVX1rV8GuG97n5lqVtCRTEOkglekYmtTVlj63rnvhE9pLZjQ0tiuNAp9szp9dU/l8SVAnLHmwpJ+Y4kojhtHL3GV
nWN17tzWfU/U2AIe1shYUaMjqWLndd2NuyBPaQf3NUTo5NV2cTYXIOKLO1kSET26uASV0O9EFGtPqbhf0uJYJXUp1SuOMh2sQEue9GtwC9vRS6GUDc8782Nxr9qGJbkV
j55S+nNoY0hl4qp9nKiNRnqbGb8TecFJ7LNnEEbJ74BIHqOfEHsLTpHSbi5HZyKygbP2jHfPwdf+jdeXa4giHTJF+D4Fibhlqs75EjZJyqQhLacic8VL07m2zvnTTFr6
9UZJLvY015YtKog8G+HhPmSNvujCRsLrRe9Ukc5bPJQ5KwIbNO6TJ21pjVK51UGfJ+3yePOgtl8mSNUQDcZSih0PO8KM1PvuLY2mOQA86bweJ5WzZD2GEpiblnhPS4ZI
672JKnqF9K0ywnGEfJXe1ZCXtHUbvcnUrHQDnnoZso7Ndd/B35OZY4A3zPCdRO3YyiLwlfMt2Yivn5shr19z0yTeDJtmu5VRlx0U7YHcu4WApjcc4q02He313LOLF1SE
WAX0aSq8jdPnfYofg3WoHWdg+vqPZwvQy3BV3uRsjtogdAy8kJ8fiE1xMrYpTQkOB9/RJjjFTJ8Sm/6AG3SccfFRO6fdNnzdw04iO/ld7NTwyZMGKvL9+243Bu1zLuCV
idtGL4/jtsQRdkvvU6gUNzs+FcowHIPWZY/nMBcBQ15fYp9T1ZGI6TxHkzm7RNvfZI2+6MJGwutF71SRzls8lHUnQ+YUme6cHLVwvBeQHXmgYzL1vb1H3RvZydSoamXi
bXB6hjooycAC+LdJgAPDHZDdT2rcUC5+gEQ/BhhH+/X8CR/2rT/82NE6FLUZfS0Ayogm0Sa9h4GMq195YwJtiDl8Po5ZijgsovSgKJoiE/Z4Ksd2jPoaqy9Kcxex+RgG
fxcLnQylypxZnRLmA93hsKxo+wc+Kb/Rqw2u2TeAZ8C7HMoXjBgX9ve/tbOcOUgjL+Sr9OKSR/nWt0s6uRxw6jxQogrHIgddBkz/1N+H8D3QhqLkVIXJR0fyDUFsj6PO
U4bUgiQm50jos+tlrrpgYjcjGH55KN2uR79TQUaBcuC5jnP9SIdSrCwe+Y6uV6lE1Q37+KyU/7b0gCx5mM0BOPvh6Uf3+WRm1wZ0zox/8chEx7SDuyF0S5IAc1wGiFcJ
j/km7jaTd/ZUSRcYQQcAweKArTogNygt1H6BoSO6EGysjFJcxtRsr8yMUfcWoBKIkN/LXRDp3/boPfCBcl+/RzCx9q3fK4LDXR9svPdXVWlrpyRfuwEkJY+YJSf6Yu93
zq4do9EdH9Ty4IxkXdXPFWRHn/75T+j2SValZgUwGqY3UzEegYSZZxkQja7FAngXX1P/Sl47oN0opsaBjYfRUjM8RKzVrX5d3ZJyb8zHQZHKhutP56KtseqsBQIPMSVz
qUFj1PB9ykGEmdKri3hgmAyKb8ztDaaGdHowT0ZJLfwiGP8sbF0njmT7/2yI8rkqRhiCCCYWJPkXgKWlJSn38MJZNVnPyVuvmFYQRFWbwwsPeffbmCYAxzf+KYgk8/dq
IR8wcMKy+hiKKHq6JXcAiu5BRqqKCWWMFvQb5FifQfRLZ8LmNOiLDSFI0TxFfgfcFnZWicTzRq9LDr4F/NM38Lwt/DWVWEsBVYsBt8WCoUlvbqY/6j+8yYy0Wg5Fuukq
Vqs5PsmLUBHURBgQiQl+4oawG0gTXycvwFk9+F4zXagiHFvSCu/TgJQHIRIKaK3kkJe0dRu9ydSsdAOeehmyjkwIYg9lPNh/wfdHfgtMSysreMsyUcDMG7T6frz2BeQR
Cg9JJGW0kkQ3L2EV3q50PfmsWvIOIKOdpnMn/JV8B8byTOgmPOBGXLUPdIaNm9J6N4bG1+FB5mRDaxhLaxOh9uWoP8tj6dXxcllMS5oJnwuTKM1u+2Wg4xOxaWGRQL5K
RhiCCCYWJPkXgKWlJSn38NIS8xbceiuex1wqpoTk8655QD1udW8RCwLIbtgfjLcx3Cd5h+guj0Q0QK00oUouaI2KPywLPBFk2uslM6yjFD0hGBZNPgV/LQrQ/F9rx2Y2
N1MxHoGEmWcZEI2uxQJ4F19T/0peO6DdKKbGgY2H0VJvOQGQcxrIWBV6sL0DADpQCgy0NKkAjaL1LnsSPycgeQoPSSRltJJENy9hFd6udD0Afaham0WzHchsil4N3FwW
96Wq8DC1lq4rVuV85fv8BDFjjywmAqxunBI6bKeIL98HZARyXv3MRI6JHQ5nGHAD3fhhj40lGPf3MwO93X/YLK040h5ouG8/9bxKZBSiRBJz4NZRGDjGg/Yxn55ks3aU
XbQUe8QmFCI+YDTLKyjSoic9TI8VVfxwqk77JJv5rcj/D0De1TVb+B2Iw+EDIi20U8Mu4sutT5OyFMUxv6aarTFiZ/1N++J5mriLX7iVoF4+HW5HWjEmwWiDxvtBc5mj
Qx6m42++mJ8oNPyoH+/Kvw09ijq7E/YI8fcKPbpp0T+sOwNdD2O7xyrwoPZsR15YirD2soG1jAoLYz/nWEtaylyNPqH07BPPZosnctPzry2IkaK4e9UE/wBZXHHmPqpN
lBa1yGo3h/SIX3pCNmAW7+00VYG8MAXhwWkS4ag+aQoomrh47GCPOWCiO8E4BHJcGZ/LQK96Rpg0/h+7SCGiucjyuFJ3ILCA8+LwgzB9orrvUEV5WwDsrYSx21rN8XKN
jtETOQpbSl0YcVEdPgA7cjjbm1L4xgG6mxVIkr2ktTK3i2idn+4+yAXWCD9twfyrxYnjRR//UucNfkhyRgw/FWTFUPwtPqLVJ5eRwjIxq+Nt8tTKrrou4j0AwEPh/h2i
R37O5y0fVhMrkdgAYADV+aI9xyiex8trs3ybmga+jSni2fdnhwfwfELETMaPFFR85vNhdV0LGYzvr1AksX8xScyPO0PjpT8b1V66OXyPwcky+VtzLVZZpxD1KAxjbZbD
Jeew59te6St251ysQfBBAfW8679FeBA3hwFLhrtpj/ZcNU9hRRl1fsVU5gLFR7L4hrAbSBNfJy/AWT34XjNdqJh2FBvIyehPz45z54UKybYX7XXCcBFe9Gpd5hJRLxGX
oZJDR/hNWH11g2gAh69kAFyHvkU0lmCRgdC1Eyk8Z3s3hsbX4UHmZENrGEtrE6H27j/+b2QfroeyrXd8KxSj+jK44Ag4yvVbzlcngQSzdP/YrenCpejawqDDUwDSiut7
DGGjYSX/mJhUZdMFPwZj1ug8I4DVAGqLGtLDlFpSh1f01RRVHzTIWO+VP4bUHWnCtFORm0LjyxxPfLlI4FPKLZDF+xfu4ZNyscJBSqfM92A/FM2llkPWADM/qhndXRiK
FlzvMALyxPsuDlcfuWxeXIX6qIqqOJW4l7fekBAk2hGCsr9x9c98JZgJM75PSugD39Wk4AhZ3BEDO4V3PggEpA5tbGcN3MaHssrwflgouCtUE6CjAtb3NS5A+9SOfXg1
RuRTR9FJ1S/Fmscm7eMKUVL1bVEYSLCZ0J/fAabV6BwTQmCXM64MqLXqAock+MHwvAVj+rTsn1XR/BYljEZDNbd/nqvaqZJxOSqeFaZAgmxc87IOTcgLSaToZt+lYHjU
w+z8k5BDj9Eh0FAsb9CUkiB0DLyQnx+ITXEytilNCQ4eUfn+3awzoy6DEogQ++XRYm7g4njev+mCxidod3fMkqr1MG9bNrQmD+ryUSecVUoeZwTMC0/rBJXC5QKs6vNw
32s95RXLSZWCZwoNJPg0/toWJInSZBymPzhpJQ96h7ZXjeksZagXn3S58X5RpPu0cD1fqi8OcQy1US/UzandQnBu9ZZdFNZIMbh6monbUE726CKMzl2KYXkzYGUqjjmq
6kp6ncrgoqvV9yseyx3W/L5ijulTHEfXaydWVDNKlisW7ec+eIYjHEbvWKvWEOemfvlpS+vpSmNu4ld+HTVI72oXrCIxHzrvEwpnRV/OyTpK8wcBwVTy3BIqW7RTCMYH
tFORm0LjyxxPfLlI4FPKLal4IREO3miLcDSiGhQaosBInWFYPFsw7EK4BKvgzqB6p1794s9IWGLfNx/bN+CFKUoBELkgTYRTKQljRiUfAoVgCnecd+6kun1o+BnpYnx+
PdLbCg07l9TH9jPvDKVKVMJiSLwI6HSo4gtLxWoN4CgzlCveq0vMQePGY8kWctn/CrM6p40+kVsQhHCWrnmBBf/CXUpk5+CNpJZ/y0JpHi/SLqvLRTcpQdsgx42J9476
sqhmQca+4YPu4ZxmDXc+qL0FWEPtS/suI3w0OR73UZfPF2QtMxaQqBhCRalJsfWefAGxopsBcL7c4aIPml8uGnZ0+GAsYscL9C4bvLwiojFVQ+4YD+qikOjYLhDAPd63
KJq4eOxgjzlgojvBOARyXDg9eDWxzcWtA4ZrPrXhiN5i2RIWkdaZQ830XyjwA3sq9tH1f3wxiT83NHM+eQUFBMXB+yrBnUiLrfPY3F756RYD0HcczqJnHi/FodaWHJEc
q1fNZUwlhQc38s3KNghadoR+qSld+IIbqqnJyrU6tuI4hy6TSSfuYe1oepUtdDS81Fn0uaRO5eThlMxxxnZmrnwBsaKbAXC+3OGiD5pfLhqGGEwyiy2MyE4t5dZAwquR
SB6jnxB7C06R0m4uR2cislq3u/7iMS9hh+auJDVAr6ysuwInihtl4Yw6afP7tpTXo21eZziZFthSrjJrcx9ZLQmMOkXoYpEqVjJ1Hm+f7+DlFmTx7QtPso9jTsLqu5ai
DGGjYSX/mJhUZdMFPwZj1rmNd1QoNj+7BMIyBTB6r4yqoHCeT9M8/pYY/S9K8kZd3md/GfD5TXBVSUpWGEOQImyp+VBCTnVLO9RT4ainGymqS0KjFViiAE5sydEI7GeR
Kvui+vmTinfHMHcjiprKfbkLFMlv7n4DS1GVQUJFu0uf/UQZnPRRF87cDK5rDArCRFrFoMMmmtr/3GM92kLFoE9+Lx9azigA9vM3sVYCu+g3hsbX4UHmZENrGEtrE6H2
clFL/z8aux3g/IAwB4e4l+cZIAameYKFXIexRzF2g9pkXzBiDeVc1PKVUASZLf4wwlP1dAPHkidooR1977U6lUraIhH7VWq4c0d0owjUU7KZvVMhTVYJ+9w9LESr7+Y7
oUQwXnDzEP7FJxljffVaqM/W+CFGmauYv7EA6L3pJctIHqOfEHsLTpHSbi5HZyKyU00B1/niPZHu0aaejPybWKHZZi+MFlQW79dVZQ57WJNBkC/ZWu25nUg22jIrKvjr
y3ybeEBT8oTAqTd17TfXUyOjGTifiVO4i6PsXVEgZRIbZtTogeky0TRLdh/Og77yesF/um1itLc2fJs+OKHzx9IS8xbceiuex1wqpoTk867ybXayBknLYY+ZHbkV4R1N
Uqywf75stI/hx9vi77dxJhaVEk5D6Ah7h51Z8c4zGV6pQWPU8H3KQYSZ0quLeGCYoyE/FLbHz1yaKaFOl3iNCQJIods6B83CNUZD9iO4qpsX0oFCyfEkr85n5fIsY15O
js4twf49qYPpj2rqyI8+BzeGxtfhQeZkQ2sYS2sTofa1jUvJZiOAjL2hHejbg+EcCYw6RehikSpWMnUeb5/v4It1oOvgL+h3nNsNU3ujf2Z1QlQP0dzJ9XRwT9HHAKyf
MAImfJQ6WhNUBI7VKDk2CAnXgAu6J9uGJLrab949aUrvE2x9KdrA+nTjXyN2og9YAOjedpyLtg1IjLnYMAfRPPRJjX+w4yoR8i8TDEBFEoPJv22KIwr5DTzyiw8bT/PM
PvZFdPEUL85OC667vhxFQCz/n5BpNajmwvzB0QADsVu1EcBRW9zltXp1JQEnapg4qUFj1PB9ykGEmdKri3hgmIanl4/BXEf2FZHcC/AnCkkCSKHbOgfNwjVGQ/YjuKqb
339lq4Dk1q6A0SpNP6tQgX2I8AmNmXBsXYUlSYNsK10t6OlvimpmP03c9FFkCcPB25jYwINSGHwaQhq2yohUJIcaRNrjJm/3cR/W8AhbUOlAEOY24sIkYsZTL8wivJJE
Ytr3oz2ykbYCD2mU3HmCsodpGRRfrRBgKkYo0Q8o1e6WTDZ0w1fqDSVNN6mfqvptlxhBREdPTS6LNg7VeEK1pJLj2ZZMOeKkXvwd0xbcmbXm9GLs8yWYbs3aOiQXweGh
FeDs+AiJv1hVXsME5i+gXpF3clOfVIMBhIpmjJJCnUnOH2FHC2/36yb+3GxaJaypenHODYJ9dIlqeBNB7M5UkKy7AieKG2XhjDpp8/u2lNdBTGp2LZiiZWT09hnlnoP3
ORfVlKXcmChrehfMCXEcQXTkBpTX52Q/OHkwyWCxAIo1/XRrESg1M8ZCxZnM7nBzzmHa2j2aRO1XJ/klG+rR36rkzd+f6QDsJZzvv++oEau4s2fJHy21cULPM8FYYomW
dOQGlNfnZD84eTDJYLEAinKELGZEpGUNlRE5YV1ecz2m2rpGoYDB3ColNfycouxN2/kCIcUfW+/KLSRTCF06Y3F5aOEJTrY4enREb7mqxT9agSCOU0gdyp5LlXXCpM4H
SB6jnxB7C06R0m4uR2cisnuGhTSMnxnv51oRnKTlprT/D0De1TVb+B2Iw+EDIi203nvqnd4Wby4RYQMl2XxEG3z5hJl7cJ5bwV1Tb9UmMvlIHqOfEHsLTpHSbi5HZyKy
UBvqQdS6NCcM+qCaTPIdnLRTkZtC48scT3y5SOBTyi1BMMfjmAwiUjDwn6W0opPfjgvPAAWX/VM0ZZ2lG3R1F0TCYqMmbE1Ia5kJjjOa56f+pQ5CjNOrsEiNKj34fv+M
CDbHeWxDyb6ZdnGu8lfRCF9T/0peO6DdKKbGgY2H0VK7vRdlYLojGRLDfVDCicCqaVPPQ01f31p6klXLonDpufxr7s2S1sDZZQKybpqrEMw3hsbX4UHmZENrGEtrE6H2
aVbbEE8xLGETyV3hmVJ4pkfUM9h6hf9RX2wpjGU+SfWK2672bU8If+5XQFz+E2TWUUwi9X6DEYOZUYh6ckB/PmXt2HJXnHcdT6HhKe7xS8XjIQpE0lO1phtrq2NFCbQe
99ZU9Id4KkYj+jnRS1WcqQrLsMZCz36IbaBJU3l1WVsDimiRlRkARqt2XyJEqiArAvWyVONswOX1YyLp7Cpk1Ugeo58QewtOkdJuLkdnIrLquiKw069D+vx2IQCOzZJa
ruTm4ki5Z7jQ33I/y/hkysB78BNz1ZALGigHk4xQ97uIiNwNFIgmCK8Z5ylQjoOOtNkE1Xbxwdl6RBye7dPKqwTmWxiJpo2vqut5pPy6FVheNxvozgXCviJlhw0NNlFp
GOVlbVt0U6ONusM4Hfn75rTZBNV28cHZekQcnu3TyquaGSj+DTKIX4nbgZNrUirvN4bG1+FB5mRDaxhLaxOh9liUnVKfG3ySEphz7CKdAl8GVm676/cFdH2Fh7/AKtjY
0lHGNsO1859rdKIIYzWjrIWBFZy2CJjDbwEl21QfW6NjuTtlEGdnyxlN4Qi4gCAm7TCjhRtjchq5YWHVl422H7OoTKgVLdV7IAH1ThUMXZiu5ObiSLlnuNDfcj/L+GTK
wHvwE3PVkAsaKAeTjFD3u2u+CBzJv8SFX2bbiAXdKAJXzpKbqZb3hnxOrDH5FhYCa15dqCjXp4HzXH2OKptljx9R3PRV5qUAmPoTNbVGAlUxbKZEDQHqsJLJkvGcWL+g
VFZ7zDqsRBu+5aSMK+mlPoK44JU5nJTALDLQunBjl7BeYhkPYPIkZ5I7JLPAbKQZqpmqWKdJ9xKIn4qYuvwJbP7YRtnE+2nJSxaZI8kfIngGvs8MkRMQkyOs3MFqjFYB
CsRdrfbG9S5T0evEJzMxN9//K4yhmN3UJuKcd3tv8f8XTc4/JEFp8z6TwHSmzfg9hD/U9e5g1dNJeDcheRT8/7O7HQclXri+0xClP+xyHToq+6L6+ZOKd8cwdyOKmsp9
RjKU8g9fsuJeFSd+WM2FhrO7HQclXri+0xClP+xyHTqty3VPRzOGP2PNeUevKxBV9x/mp4ApxSnoHTfdx3LhH7iqaRIDuuEKVcdSm224n+llQ9vLw77LrvK2xMxv0gfB
sY8/i+QR5m0XQhtbWigXdV4vQ8Al+RH5+ASpotl/QY5qBR17tWQpht24Vd8GxHAhzYb2cwqjlQcdinRrs9LUTsMBUSLi3Sc6sR7Ti6N7EWe4qmkSA7rhClXHUpttuJ/p
SEE/RIUPM/uKy+F7A5BNIeWj6nh4216pAuFcOfF/WWE3NUnfiyty03DlhphZok9lkP2Bg6tjhRPDmKTS1tSsnA7f6diZ6LcPrbzrI1dj4T1wq6thrXN0ZeMdX0aEeFr5
sRQ+RDxXwUZdXFf0oaK5m9ZtoZBUsexXJ/XsjzYh6ZKjApTHGKZZBWEaq+fwv3mnWjbPvEqqHqFae1afe3QVAqWZZCM3zHT43v4JSj4qBVbEflZXzMFOBSQx9LpXCgAS
Y7puGkkhvKrgqiSX8WQUm0DM/mbbvp9wVwvxHJr9WXz2BWplTn7jIXOuORfkjeZnTdgNr/dB4wlAG6iUulQJ/gU9xzAQS+n0r5a2USIkY4v1Um+mU4o4Wbx/6+WNjiYm
I71ucW9n4zR4xTBpXuwvaw6DYokudE7EWxIVWdGNZNz7Kd1DqX39x8sC/tFjflrleoI3KRhUOSk8cwe/YuUC8ZE4icis5OrQk9tI65gbiVJjum4aSSG8quCqJJfxZBSb
3HQK4rxiyZQhwUse1FYuPTJgobfkGY9dVEmZoIvwirG73vPPdCnHtPCGUOaE5dm3+XDNjhQoIo4ApkRyNHCOYGvxBwNpuJJigMjNh/HBNyf5tKsfn+fNnnQFKLvRq8BW
fo4caM0NmPzUCZPHluPwZBDAOfznDwkSHiWrzRhS+lWfAknoNGvtQjT44rd7iCoxNDKHTj7KtaZG6qws6/3Gx+SRHZ+Hu2wUSu5F3uyuI4bXT4ohewVhM4bpvRq63Zq3
FvfYB2g9F0uklOC5xS1etOTFaXqtmtj/AImGbolcQaq8FtBg1+VwaYpiwU31QRn0WacfroFni2ABS3NE4SdwRmBeJDFK6t0ksyb5UF2l6fgKD0kkZbSSRDcvYRXernQ9
v3iw46Vp+YrHHw/jYh/ld5ouq9vSxfsdtqT9AhODhBgyX/1jCZ3Hs5RBdN+jccmf7kFGqooJZYwW9BvkWJ9B9NVgPTCsLiLTz6cQxq3Ukc9HVj2/YgybPTyxNFVxspNN
vwzdEaOWJI3ms08TKjHOuhoYHbIWLpA4x6jtcndmW6Y76izWqSxCIHy3gEbUQnwqNrdMQwYWxtBVgdzW9+lBIRmIpx3pIfrya2JeI3X9aGpz4iyUqOsVyRTtaBR6YvBL
anz2pT/yYWzRDwYoQOeWDIj+41bml+OhWPwdisz+wZqho7kR3OxALiPCEkkprpMDs6hMqBUt1XsgAfVOFQxdmGZtXdzAtyTo1J3/B+b1/rG5N3aaZpJT4eptC2UFnOdf
fcm2hG+IOPXPFN/6VeGMmc0bztDHoUw06ZVI+C++HZRjo12PLbVN7KVDSIWuqNueAcTvF8gwooMKmKArv5m08M1NQtkMovcEpjB8F5S4R1dISMtDGVasjdu5SfDKcJqw
zI87Q+OlPxvVXro5fI/BybbjmmsHloTdsIHxLTq3giD8CvFL9nXrqXZvAioIb0/7qUFj1PB9ykGEmdKri3hgmMCAc63vb1qKWNRUIePOowVAEOY24sIkYsZTL8wivJJE
079otScYjbwOr9FdePuu/QHE7xfIMKKDCpigK7+ZtPA0hv90GjHKmVIv4cwwdwHcQxRRcTHR/+ipyxKIJx40tc1D9qrbkEyUFah3sU9tLUf2jrwXWZGBN7DpGIm0ac2e
N4bG1+FB5mRDaxhLaxOh9sY1kqBQRus1x/0MghJoNARgIyOtvH446IYNRReECm23lM9LFDk5XemfePQjdp0FiHdQI/5vW3pAEDtJ7UoGPAOSBNyx2r0dBxrGU3SnHfzD
swfBMdQa9YuxFQ7XUOdxABB9JNhCSDvpMMis+OzcLLL2jrwXWZGBN7DpGIm0ac2eN4bG1+FB5mRDaxhLaxOh9pXw+NSqYOz/XeNya3PPRwUzlCveq0vMQePGY8kWctn/
lnzk6ZfKnOh88bUMeIxU8pTPSxQ5OV3pn3j0I3adBYjIBAhwAjRGaWTsCwtemgqsU9q3nWGe3+BUuk6qZ7Ydhh1nvnIpgiOC6AMbjj/rccbMz0Blz1sziQU5Z4CVtMMK
YB52PVJMTR9tE+5/4tgs+FK17gpyqVKvGWdXgA+b5syUEZ/0bWguMC0dZ04NCWTnnSSqVw8/wHqSonyLA9/sWJgAS//CDF9OepWJUNzoGTWjP2KDJLCZ2aGToRU61FZp
kjJnbzPMZXiS5WtN19CASyVoocTCXU2t8ieP9v+j6lXMz0Blz1sziQU5Z4CVtMMKYB52PVJMTR9tE+5/4tgs+APknTgfOnf1r2VVMuu1RDTLum6X9JKMqRIWmkykCsmc
QmvW74fUH4SNshZ9WsMWnZ0kqlcPP8B6kqJ8iwPf7FgVjoG92xmURnHy+7JLYLFXcCWvdTJftzThLcocwdCKvJIpInE4sY3vp4ij8wPIStzRJ5WcMuB+Z7UMW3x+dWE0
vwzdEaOWJI3ms08TKjHOuhoYHbIWLpA4x6jtcndmW6Yom1bG3inHat5v+ZbCDduoK7eKeCXPW9LayrVc0CXxFM0tWuONOKZGTPPdpRHyekpKnxyyElTNAM+c0BRAgdO6
n4Gt8+8X7V2RYSIQ3e2IZ1PPSxBcfcxVu1XdxnPQeUoBL9ZFQcZPPqoW64PdBVNbM3I4hMF1gAZsE5Rz2X02K+Y9wofYoU0er6HUrtwhnRqqZgf1Sru0vgMtJIeqEpMb
ol9b4BpyvukZDRA5O59XK9h9DEmmf8SwWgh0ZB0+gLBI2mXNuGkksdCPxqUqQZRMW8tmuNXwU92bqoFW5eDGdwl+b/TixI4Ikx6Qn4ywrzvmvf6vlELHdYiUAfkPEJEu
StoiEftVarhzR3SjCNRTsgjs8vtlbyNfYj2sNd/5t2OKbydLh8XThvegMKG/afjo0X+gntjanA5WTo4klhgV4VWSV3m0i4z6B5KS/yq1JD87oeBURpzihLXJC+iSlM7a
N4bG1+FB5mRDaxhLaxOh9s/iToBK1QzBSLHHkrriboczlCveq0vMQePGY8kWctn/gVqO0oRX/MDo+qwxWX4B2UQJ9l+iZaG1h6EktoXqwX3/e9DDKnwyK3q8A1s7U4Wm
qUFj1PB9ykGEmdKri3hgmL/1nugWN/9ih5iVKhZ28bNAEOY24sIkYsZTL8wivJJEYtr3oz2ykbYCD2mU3HmCsi5QQCmc3p0IayDMcrKXkQ+FS06zdohVLBPFMm3NGe+f
Cg9JJGW0kkQ3L2EV3q50PYS0T6EOKTiWuNDPDROmOboHPZWQsl53sWMdpIBYDzhjcHFrY/rzrbziFoHfpoRppWxwA7o3gvGYX0l1sQ+2FODLv2UQzZlDarKkzEDIZz0b
aRBEtvy6MXh0X5U1F3+XSuqE40m7n2X7dejjOC9fsAH15ZJMlj++VnlA5L+pKGRr04whBKcIehW8/C0YNG+CGodGE179D8Imr2knTM+eQi0jxn9mPR3kIrLqA0qhIwsj
aa7Yof3LZaYMsl/3v+1TahZLBAUq8f0pV6cXGy7cYJykBoyZb44ggGmmKtC1+rL+64dtjMV27BHi7fwhMykDO47XVL0ze9KBxGHhzoIbtSPon/ef4WLI7JJ7+ExxnP60
a/l3j5n1TYLZvc3E+HJmAGuOQEBPgr0W7RC39cz56aIPhNnN5ZY7aUUSwrM1m3FNUOFJwZAyKwEwZu7HtI6lfLipdSo/aOPVGl8a9c7UCRxdRokC9Xhw5jNpwDHa3JWe
2suyFT0OyDthqmJaAr2uKWvTc9Z2Q7TTu0dfuaEwHY2WJTMrjDUhV8Yy6ShBIjcBudCCyT7mifMYsYmKvNUekOAtjm9fBTXu7oDyIowsBTpYBfRpKryN0+d9ih+Ddagd
Cjea9F7BbcCJN2cyxT+jD8sovmS2rKcfJcZLE8rN9vVYBfRpKryN0+d9ih+Ddagdh9WirKh4/pEILI5m0ZG0aBJkIZAg9NEilk2WnQuHesZIBEL7VufQBhr4V558HR73
rddmiMEmRm7HLkdo7moRzzUyRe71xG4CNEQk+ozEGuGRKV+PQj+FqgUS7JAAGi0kOHEXpDUYnvEfK2C9z3ASn0u2sWbsxBETtpURt7lJC+HS39wPAxTAkKHH5V/BN+gf
FrqkgyE0thwEU7ljKuYFI0IJ1QnU5UjxtySqErtRg3ge8TAkIeHvsJg2vu/BwVsC3pjliHrpPXHESNW54whttUa+SY2uk/ndwbWO7w9gcxCgXZasQWUPvZMsR/cf1fCs
QDsnC8eNBMsy7UaQJPnLfPCDqhdwxZnu//leBvYUT4NUgEDV+OVIaTgiXf2q9WLnAqp2TWW802zWcOUeiIxXra9Z+wqtCWkchuvDpukps/JGiMCQUvYgZGi6MXsDDK1e
M5xEem2TqK2cIC0m/9D/f2uOQEBPgr0W7RC39cz56aI0slkzNUmNdg//0ws45uCIxJgT0pNCgmeSk1QS4wGXgUCw+SynvTwdCFQhjT8PO/WJqbP4yNIqeyr4hoybAI97
IlWJnguEovWVZNztjgwbr+bsfNqIpQM2d2TTJhLlBGt4gjidJ7McMlVmarOUA0lGUseiV5sNdsiV3Gc/myEE1fQvUWpWPkJl3BnmoXrrR+/a2mv+SJ+Mxd9z/P1YTFPX
av6thc6grLplR1PDfqvQg1RLUwa2rymkJ1KB8TuoRHDgpTylGJBiRjb2EjcXt0yUx+unz3Ks4wA7fmHw4RYrXCxkKs4Ko4NhVUEA4Vi8kqrEmBPSk0KCZ5KTVBLjAZeB
zDEbIgQJUe++joon9NTdJ5LdM3KE93bNdXms/5ZKuOOwv6XmLGaU/dbkr6ra9uJnj2ouzgz4UN54HcG5SeH4GaM/HZ0fZnTE6qH967WUH5LLTQKawyhWTq0qzQZ12mUb
YV6Qf9vBGgEN6Q0N2dzSYSPVM+A+MgZVzOrpkdduAK9tSaPK7KmLrwyxNrV0IZnBNR/MzNbjumL21INUdvKPUdXQ9W/VSDcRv00v5kQywo3RHyG1itkklm+JfBQZSe1S
bl4xPg643ANnn3EmekRHoRCJLOS+HkbD+vejgUAUYcHq4i4yRSW/s0rNud/sgXLlMKyLFiRwqX7eVsmsMDCrmp1jde7c1n1P1NgCHtbIWFHN9v0sRC4p7fvKZSpq6MlB
KEiOABR8/Dfe2gwz2G5g5IAVFwoUFuI5PVf+NIlC2I2h+muFgtIURAqMNNR5Bdf72RSRGFSm7XHFhiZdlmAk7etepr/qhGfEhHC33IZRoRPGxFgXN0fh5ZqLrnXtEMlq
G50xSk68S+Jf6kO82xsWSZS3Se/7fBzmLnLAhx08H2sdDzvCjNT77i2NpjkAPOm88TJACquivadSPetcg5sAjjKwnbkZM8pay7kqDDnI4Kfx04JwRcQ65fLmfzZkXYaN
PTb4bmBcd5lMtSNG36CzfLAWiyIcX72Hptc56jaCNZ6wvBwE7Cmj2w/6i11JenYAXEGOIaSlpXG8hB8zF9caxu54Ad/rviiFv4GLVv7wIf548hoeZh2cPYhblve2jWO4
4TdJHCYKMSWpsA8yfj1XWLEX1WsGHTf/DURp7xfsdwXcC7xQHGH4vg4OTLIf1GpyYVhL39P6dNIiPChkpRZQ7D8/rPsW6AYhAVpUvWykTAE4rJ9PfFjqBAr0dBJrWC8E
RKtQtfm+6jCvHrfsszAwO25Tsjthtj/gbwosjjj649zmjYZGTPpx5fHkDH12aeTGq7OtzGL+nEsQfaoHtpD9HZ/Cp5FViS0iU+6DKldMfx3m8UYhoo/lwxp2GL+KAEde
eacMNP/QM4xuSPdHwr9/kYY67Ty//MtEzgKc82tGahX02XR7cVZNtCsjfPp9+JLByogm0Sa9h4GMq195YwJtiGXUvqD1Ijud4Fwsp9Nu/KIeZwTMC0/rBJXC5QKs6vNw
yT1q+LZpG0OKpQiPVSBkxfaziiK0Y7H4bep32Rr0YddpkQpKAJfcztHRAqzoAFM0Hi2Fm3Qlb3U0VoE5Fs3EyinDaoQriLhO638W+fsM/4UCTVH4MGfQE+oExg55IJRJ
rdfMEZNdgPp/L7BdyXnGxrEX1WsGHTf/DURp7xfsdwXrLQkiEU6/9bQETXvxoY3pNjbwYi3FGdv/5OLTLeGDpNU1jNLCBwiQoQRlhuekyF/hPMfiNU5F4zo1HJLP0lxG
sRfVawYdN/8NRGnvF+x3BQP1vqIF2Y9K4B+1Ga6ggmIWel5wngwbQiDd4YtXFZ8J+lK9LaN50ESehQ4hmSRjLZrOex3QGcGvrNoVlSq/BJuPZ42TjVIRYyJJ5wVspFM5
rZY+XdSkH4lY6omSSWNTV26Ocg6EJ2cM82rSSgc3XtfMB+9cadiOnkTQ0lTocvF60FivrvCLnGLHeDBtfnY2MHSkRXWW5EN/fh9WHrVOHkV0kpa3m2N5ElaiCxnBJtQn
7ByneoACUSRFLQOXVrjB/Y0Vk8xeiKdLLWp3xAJM3PA0NC1GASKTA0gH57Jb09jRkJvpXb5lkkq4GKrK/bQJs77dioBEDdM2Dl9SIooxVQ2xpwgnN+kNvLfZz1h1gfDO
TvbyRR5nuyKf2hYshUW+Uy1XAXMM3eZQNDIMd2qGeKNpkQpKAJfcztHRAqzoAFM0tSmDwxykXQkz2bW7uqkOxcy8RWTJW7KiisSsD6uE/F4By/YWj6jcVSnvfUybWU5K
MJfaHs7uaTHs8Al9KKSw0oDsxLkTm/jwvVBbwjDgflve2DfolkiNM3wPtVD1H9WyjSSZBoriwiibT9fDabDJGx5nBMwLT+sElcLlAqzq83AABoBbfY4/KhUI53DBviYj
F8rgRmL1Bm5mQAr8SKSInUdsTxHSMe8UaREA9s/I8YEFCv6HAHhNlddwZAuxc1/ssTXZlD8MbYWBbqrPOajte1mhc8hffZKXjwW1lTza2xLnS7zec7N8NlEguv84tvOZ
KsU/sOkTInMGJ3V2ccXX7uOTscoxQ9LA3IIPZ7Ge3x5de4Q+HgG1VYpo+wFUgnLK4TRkrLbTE+SXLCclIn9UVq5DK2BQ2Ah2svUArQiAmMAU9EHPTFsx9Rzf1vmGMqNp
EoGq7zwPAdQhzZfxM58JvzX6GszZfS6juBt7qYERdugCmlC1LCxW9hpGfNpxmOAIgOJG41aD5Qm+QmYnd7sO66naAyYC+br8/iSSsRCvCJC7lhQ0vJwyULlby+mDouMR
XigqrlYXT4iq8r1sqpdO+rrZabOv7PFQRZN/PrqrtNMafPzBLzGdddunS+ZUvGKucA1SSnkZ+kwuhFR2wm6V0iQQbTul7aAKL9CN6RZ7n2bnzbw/diVT/UF9Wd21e+sI
29ku/QIU11oDDkUGYBBBa8bHSE+gtaIWkJ8qXRflZaynR67k5QWltAWpj5ntd4cRzzx0K4Rj/u8sKf3q/ZjXfmvTc9Z2Q7TTu0dfuaEwHY3tXKNIshULVloRRWMcl/3Q
TxSvGMDe/sdFNQ25lop/Uiwz09FsBtkXKjZ/QniwTII6+4qH98LHP9mmENFnFHWkUvVM7pyfVT1twXrGUDL7CwfJUWQaHgbFmYkzumy43DJgsG4e6ywWR5VOJsXYrMY+
6+PqlF9kFRc0e9hRZ3/LckV1lpkq44C9MIZuh2umpQiby3AaygTfu2WmhpVgAypeUr1Wk4pGIQkks31q/iHw5UPbqN0QDnow+8j5BayNcGVTJiPI94niD6nVzmGh6yFD
1EZmFD40ajXoRQDlIbzO5mo9jS41TyOr+RxrBwPdrRRzlXJJN0SVZD767fMg1GusivlveaNNV84pj3UUY78XbN8WoGYG+2l4liGoFv30HmfPT+Z67Is3VtrEdJ/wQ/Hg
GBM6V+al23MKjaJOHQhm0NZyvMGkgPZUCXuUNpxhK5xq54fwwfDK+7UtpntXHRjWJ1roFGS2Db3OVKgpAnhmH8qIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17
L8q7MnRNTN/jkwcw82rga8qIJtEmvYeBjKtfeWMCbYia5Af2OrbDHMJ9EpAFgOGxMs6Yp83sbEijSPVFltsRMJ5DxCzEkASNymFUZ4DxMUYtJY9QZoLVtNPOjCt9XGfa
kREuwLUiVZEZ3VzbMt4M9p3uOwBJwVD7uk9dc5ViOBNIfJLwI30qbKjuXz685Hs/2oRyWKk0HGc9kFJ1BBrZD85iht8pNry23J7HGLOOydy+jJYGkLEjBeMp2ApJgYa0
BoMiHPw5GySYp51IAbs4wZ5DxCzEkASNymFUZ4DxMUajARESEEvORidmZR9x8qUSkHAhZcn7Fx467oJVunPtbTm9Lc66zmvw3hphF8yJlBB+yGZrmBneblZRmw9FMfTX
xFCLbieP94jfM3WwernLigu4ulFrZJ8GOY/zyyJZ3Wf1z1KHfHgAQ8Eusjr3kjdBdhzi+RFQjsr+3WYC+b26V8qIJtEmvYeBjKtfeWMCbYgfkvpF7mOJ/aFMeRR8SAV5
yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUZtzsUyX2oCBJNOmc+MZsVlyogm0Sa9h4GMq195YwJtiORt3OZVUTG7gUiKejQ6rAUyzpinzexsSKNI9UWW2xEw
nkPELMSQBI3KYVRngPExRi0lj1BmgtW0086MK31cZ9rKiCbRJr2HgYyrX3ljAm2Iyu3EDuo9KkrhcwA+NC0ta2FYS9/T+nTSIjwoZKUWUOxqLPE7e9hKp6QKlaCQyOJ5
RvNLUWgVRSDyLaqmkMOhGFsaFcYg3N9S8Zaz8NgiGV+HQ9MqK6uzikUAZxLt0SKZyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+9telntkUjeb0MHJS6Uu/y6
rWp0OUF9NoTt/8ALWSc96sqIJtEmvYeBjKtfeWMCbYh5hpF3lQm+EBMlGqoJ56vTQ+w01OJJfKh1N5LQB6682MvUg/lpePX5/VghbrtUw3PFW+2rwx0LrqGauMVmKpty
EDrKauVyOeU8+13wOug5vMx98/BaYDI0AY90Zr9cgeNAAcRy5TESiqh0PJAHk7ithw6QUNhifXaS5isT2i7JkNA0ukO1qf2EwrhYp+jLCx0SrPEs7473g1AqVt69heqb
Q+33v3dR7rrPB+ZL5PHGqeTzTbS6oGxkT5zMfn6cdzjhR59tWQTl1cjjQgNgG9fcjIV1ndt7/ovkBqAlzT1dTKC8Z4OMhK8mwUyzKfTeVrJF9ScvLvWwxGhT6aedwNMD
ONdC+WevDhM2+RWdriJhfQz6BrRPUzpjbmEwftKsb9XACjCrgidF+Nk31mRbhVlHzA+BAze7vM+g6uspa5HVCPs/1NRVSVylYp3Kd4GA93EUwEoefgNwuIgF4vw2hklg
RZiBpxMvEqYfuvM/2RUfsZ/VqFjCnxlhXdoRZD3jU0Gi3S3ZRrbSsoy3GXYGxxoKCnJ7gV1zUGUOfH8qL7HIr2qGbM6LUmw7f6qHnue7FkKIR7Ulzh8vncvLMHAt3ONj
MZCaO0LavKrN9Qx51u2eX68LpWdQY6af7hFgkrYYS86tJHg3VhcIqwnTKjYlVb7cmWm6f00KCk0rqMqfl+1x5RnRuy0ALrNUkv9KApqI/i5PydlR2THkv6WsTm5q/UI+
oiguVRjtw0YFOwj1UmCRN8Go9q48o3y1Xm/zfBLQ+TekWvuImD1/WjQf1aED7cNBg9Zt2FXqHDsgls4F6WU37o+wr/A3jlNuxUg1Hlss3GLYfM8hbQyFYSBPUWV6NAdC
YnH9Yw1qDfg79q51PYXTZMh/sokc8BM60UmMPf/bNHyiw+Kj3maRzlv5AVbSyi+lzD4ZPSN+bogxcp70YmdtQ9y0GpPiC3RHTuqKOAatmxTqwDGF+0IFOWoEURXIqrZ+
Xxw4g+MS5hElzPaUV+IySheav3+S2gYpr6PzSHPDMto3unmBkYhPsmbqE8qxYzkaFu6G4XHjf9bUgCXkh3XYkjx2nH+lZKqYYz0ck7z/lQe78Tk7k22zoWZ46hooHGn2
K8YzzkdApscnFbhXfbA3HFyfMdgk1zrwe8XT93htztiENe3Sxn389ZOwhpRaYzjFkHJTtNSxFxcleb8/P1siyFICkMwVgQR0AWPUy58IO/W1MXLkVlNUQ8R7RPKmDM/y
XNbdUT/S4sNSaRoTLsU/1gIJg5Xgl8bQgRq1MARkPEbaK2tqHIvVAxP2RjllXuX+8BH2yGyE2vPdwLRbUvNnatrllHtVd9S/oBxY8A9/Ouz9d2dNvYFr3wCTbuMG1Ttp
QDvN6rkZCCEOiSs2EoDxc/Ve2PwR6p/uyno8/xm1lLjDuugIyIaYxzYlgxmrZDh8FW85qGNTAQFxYaOe28RuMJullnqvk3p/pAoBEh5/7D3Mr9LkuGIG8Adzhf8rdLmJ
0ReS5XImT0+M0Z9SGH8Z67ph3CtEfmHwPnmQt8wymzry/YYYTZaOixSWCOedItccATcawxhtvi0gZYLsVr2XYnT4RUb1sfzm1lFnsQ2JYsdw9/FA0tKVJhW/uJ80tDme
VqYmR3n7UqFhCoL2EEpLAvfaxi4zU8vP1KioV7vD+aedKE7eyVuplZGgCkewwJc9FUqKvfnxvgfE7QXpEnQigTUfzMzW47pi9tSDVHbyj1HxE8qag3xOAtLGqY8PfMma
zOpDYjrkRAw42qWtbiZVhcWaTO22JZDjz68xCDOBOAvfz6bxRPR+fcZLhc00GIWnah/PyEji/qIeBj+UGyk3Cv4orRtU/7UtGVGEKZB252vObfnakk7O7mGtOXpYbAix
HJPABtTewKj3/PBZ+OprIYUmjdsauLH9Jtf3jREL6/kZHJJRbJLPYAjLg11P5QSq/ZUDL4oZXANoKsWuFnGYyzFCVxXSSE5wGptHcCWzOFg4NEQJNfwPeTyXn+mP0XQY
/NihcKmii7oo58AKcnnfRSHsmXnztDLAT1ghMWmOme5b6XdTooQwcAmMt7M9a1xoZ6laWnx0FMgByOGAFf0rERuw605c49Y94S1gLx3MM7OXvRKPouiPJ90jch1bU5oD
3UkgA7nuzWBg7ynTKL+fsZnm+GNgH7vtvlcKQxiAngUPcNmnIJ4yzpwaweVOEdpVz6JLOVfst9GZb/MNXTp2aIQFKIv2k8vK0n+Sje9hmJ93D97sQvJCrHc32ps9YFy+
Hd9xD5nRoa7goHgtT69a3DNczMiLAp4cvuzUnLmaqOQpy/54x+eJg+syIx19t1YM6+BWgyhitxYV/9HdSfQTNgo6Zhdr/xEhl0psyKdzWf0qcmlj00g0EG7k7Z6YD0Sq
YzCHrcpizycdBbBDo/5Sbv6hWBQV/EPkYu8Mmys56s62/GCQprXU7/jPtnfSygkwwhB/CPXdIz2kV71SC4Oy/UvhbY7RSZF4Nz1WQY5kQpWogSQ4fbq1Jvd16HzQuw1Q
J5GfC3ZnZE7zzPO6kPLf79h9DEmmf8SwWgh0ZB0+gLCkcJNjB2D2K8TukJX2kNMkPifFznQ+SuBdgStlL2zANf/f0lscVhlnWnIUQf+6U6JSYkenNAZtOMrbZWlwvBNd
ig7p7+ZMRHhCzvpk9eSSLnDRschddASvTc7zlBpw66+kBR6MrbqsieYWviDOinCLDG7FMn6vROzsu51gtvI7XdOyxFPawwikuWmPLmdTBK192O16zljRPOwLh9QF9ise
PbQJ8zI2c7LHXlbsfbwnLcVOn/SlqpQqUXfksPxXuUWRCFafSqUOwyA44/qu1yYSuGWuIjhi8JrAJNttKAit6aQtlgvq5Hp/YwOX8NE5+nnPtt9EMKhmLPumw2ztqJxa
2/bKtlshAIdjfLyduhFtRr7vdQzU87ZUo7EKDz49SYE/fIQfsoBlbqoLi1LXZ9Ctaiz1PHQ9ssl3lrD+2Jtvmfa4ziBXSKCpe4VyfQrDEERwO1hbbWDVREueQDInwxTZ
ZRPyKU4gaHjSnS5UYLSYBWrjWIUKEC/pwvlwLzu9CgYM/WymFXJi/if3lKTpinc4unN5S9AEiOPsa64q5IVNtsSjGhk0kiu7BdUT2PrLq+C0iHIiCEXxPQtEpptUQILy
RYZ7NPfQGbc6OCgxqHdiplK3BJgpWT/bhvqrFVsWdpsXz2xB9BHQuCZiw+BNkAJoKBKzX4TSp8HIWyQeY8lGuhjbB4x6xHE/qfcQjTqd0hZJQoy0zi6OCyL6l495VScY
moRGZNRfaYx2oBK+jdriyyoE0mCItbxFBCy54RJ0XS0bW6HmTSzpHTlAqycEo6AAs+rOB76DbYGn50lpAm8GwKjRaadY9ro4fUkz/zxQzEUoWmQvh3+bz7EhqdUf9fxx
hJLhOOB+JXt+WwM5+3oMm7pzeUvQBIjj7GuuKuSFTbY4e/kZpkmyrLDPXNy0Cqfs2eJ9Dk9Lqwj2JbClOgbKWtDzsoPuphWkPxrx2BE57dom8gqgDX/QQI2YwiORqshu
lzMecSd67Rmuo6sBk007rx++HnzKPbOV/cbUOlG7AeEuYpGIjaUi7tf3s84xauPrvLG51KmypZRr/TbD5M1OZlDhScGQMisBMGbux7SOpXx552et238vJqaJkbGMsJgF
N3rFS/MhVr+8jp8v9//W6uO1HvdGPoP4dMYCtIC2S+POoyap1ey97nKUyDMHh4Vsx+Ok/veV2Bo+IS7FXO5rZR7xMCQh4e+wmDa+78HBWwLOoyap1ey97nKUyDMHh4Vs
bjFWSJsOIS68puVL4ooWgrb1aRqCVh50WBDzhlIeqeWfOnPSf0vWvLF8bzh8yTrNzuefEmoLmFZRRnrOy9SiZVFOwyhTx5cDOTXF4MtRC5bOoyap1ey97nKUyDMHh4Vs
/ugmZjgqVjzhpUvDz/mexqH7teqKoMtB0nAEA/UixGuGP/XBvfU7mbXfpicFvSPpKD5HOWhe3VLZnvwDShPjwR7bMSAVSILOJZswQ3IGStmGP/XBvfU7mbXfpicFvSPp
Wza8tg2OcMzQsJodn6msHvmJBPFab9sxTnVJR1xte+vOoyap1ey97nKUyDMHh4VsQgnVCdTlSPG3JKoSu1GDeB7xMCQh4e+wmDa+78HBWwLOoyap1ey97nKUyDMHh4Vs
hKvHl891MY3g/eYWPeVCwOXViEHhbuAwiyU1Wo31MLs+skKtEu8Q9qq2ogzA/+PFMvgs2hFDhe1xCytFpbVWZW1GRFDKQqbqBO/Mq+BRLeTOoyap1ey97nKUyDMHh4Vs
wie87lGu7xV7xxbrCrB8/GuOQEBPgr0W7RC39cz56aLnpr4bCXOKyOfoxiA0SZZF6Q8BBGb8j46oeCkjVW0gqJCXtHUbvcnUrHQDnnoZso7oEH1mAz62Xart8BPlreyg
K3LAg/8tfQCC2K7s7gi0J0VE1+knB7LqxrTiFza4jEKiD2i7h6VtdKvwvNuwisdtqA95FKKKIFIus0zov+gm9ruyOtYoZFv1muWIwq/6OkiwZ9A7BKjb8m+nOc9m5s4q
HvEwJCHh77CYNr7vwcFbAl6k0uLZI23lK3OXOsPWB1ckaaaSxkgd+F0e6zuL381ozO6mtCuj8ZJjH9KRWzF8pbuyOtYoZFv1muWIwq/6OkgcZGvj1GyajnneO8TJFTFb
B1DsRF/Tx2Hu3FlQHzO5NzVS/74WcbeOoWx+tCgrLD+g+PdfC/mxgZV7kRssJ1xvvHjA1N5MKvBegLAs/vkGczVS/74WcbeOoWx+tCgrLD9LtrFm7MQRE7aVEbe5SQvh
0t/cDwMUwJChx+VfwTfoH7uyOtYoZFv1muWIwq/6OkiiyMGDnNG/fZSWNS0sGviKqA95FKKKIFIus0zov+gm9ruyOtYoZFv1muWIwq/6OkiIIzWTK++Xc7nN2nGSlOYr
kuuhhq4mVW1kDGh6tUBNx8YxbeozPejBJ4gDsuqOHR7ftTvS5k8jzHXWUNfjgyprLn2d2Ok9xoyrq4KhlSBP0ruyOtYoZFv1muWIwq/6OkjIyYhPf6F5ZpGvtSopBmku
fphmSvaqgov8aJB+sQ3X/fYEdGX/h4V593SaL5hBxbepW7oydoEIzKy5bz5sXfa0kJe0dRu9ydSsdAOeehmyjqhd5Xztd8GtZ2gEjroLxO3V4sLom+G23LtYl9EzE/5k
qPm/1ECJU0wvTWgj1Ei2H8SYE9KTQoJnkpNUEuMBl4E8nNYXyqVPZqEFf4XvIdWzlmTBv/Jsyh2wrXC7dMiOomu+Z8LRtK1kpeatUaGlilifdmAxPf3RUk4JxFuSjN/V
/34jCL9I+3pV518U5MJrYpz2JNPCPPTythgTLdgYSzRQ4UnBkDIrATBm7se0jqV8IsvDEyu1b2gMeluIeSJ/ZjuSNr4hZRtpn1cdKDxkn3MYXOTxVuYCe9EBh9SQjfY7
8GI2KSROq+ucj/sD+faBdLC/peYsZpT91uSvqtr24mciYjAN4sjdzVGthQYzOg3goT7ituswypICO+DwQ2GE0Wu+Z8LRtK1kpeatUaGlilhL0aRLzytnIILdAPt7Kkjm
y00CmsMoVk6tKs0GddplG3AgObiD1Y6Q8DyTeAckaGDEmBPSk0KCZ5KTVBLjAZeB+DDMf3bInXJj3pmztFbtBFikODnSsLc7IO9heUAqKrDhpXZM76jFmmH61BlArXAx
ByPiqAWiX2iQp1luT0JbIBVDvPo3t+z2u0XO9fNVtsCp1Gj2PKJHeJoKlw8hLzLs+J9h+KovGBMCYQa/Mj5O99mJHxwYL95xIqnL7VIOKIxYBfRpKryN0+d9ih+Ddagd
y+/KBcRvy6e+qn/l5K8lCnisrhXNh6j+0GMeCIT5fuUKQNYwlijrpw1EVk7s170YY7ax05j2ISuDlExTeWhe1kkjZ8BXjEBfqiWydmcDiOywz6ws4LfIaOjE8aAGj72J
xw4E3kbv1NDlo7UYp1NazIuSKXRQnA/hVU287DW/ftnzXKFbX1Ptk0oJlTLTHLhIgYEsXK3n47fHF/xXpmDOs0Ja5AWAw+HlPRg32f3j4NRcdUp4KMORFMWLS6DklqwH
R2xPEdIx7xRpEQD2z8jxgYOm7KboRKxSsb83NVlHFb5DG8FYtsToNw+ZZH2gkWrcs6NCDA6CVvp9NeUYaPqp5DHjWOp/b6pH7pfDaIuJ6yZ8eDR2xoW//8E5wOIljPT7
gC3u3ozCFAcJgj5iA6NGSaWdT/FY0IkPzGAABRqJbPrpcSX2gHMBPhbB9+/QKE+PUoaSB4PwCKWe1YVCe4ZMN6M+QEpGsU94h5kPYh6ekMre2DfolkiNM3wPtVD1H9Wy
xiHNXi5uSHZdjsYo1PBF2ChUcgoxtL5qmxVnrMJ7+6bfTGQmVTAc1WWBgJa/S+BhflMC5EmLGrwW1HuZZmlKNjlCf+SKQmwiO73cVfez6pJeE7KcA9RmoNscYLwsZdyr
IOG4W1aFTUfJefrZofanFmdWjGi78idoW9uXhbVLjT/MB+9cadiOnkTQ0lTocvF6dk2lyapJHZHpSrp2MumNsX41kE++S/08ikhQh6eDx3BHrCRYTYNfvzqfJo5dCohc
ncKozQKYhnXcVRmbqNNwdlWJ0jdMg1ZtoWNA6poz4SI60tRa1KMw2akhZHuMEcXy37Dy6ALDa869V+CnksHtmWAb3UexiBcHcC8MOHt5fE/Rrv2ROASh/YFy67kPGKn+
SxKBipoPfWqAZeEUjJuWyCoubnPhoGxmL7QrRFJsJycUIEjmifdakKYyd4YkfXrEzmrUQUA/9cOxiEuh/M6uoeWWhx5La+HdUHo/vRiLX/vveX6r13P5Okg/Ddcy6vxp
O2boA1ypWpLi51OWrwkRwc5q1EFAP/XDsYhLofzOrqEnVZVtrZP9+vTNTB3QvZ0p6Dq2P4esNgd/OEYAqCH8eBRA70+IoDko9FAuBywEDXk6ymPqAQYMStftXN8c/n7Z
zrJQvcfBLZ8iY32ldFXeF64A0FhBhVPrChKkmUv77uHwHJMK8r1p9Ufw0ZnU1MbwfLCbZJZx5xvRZmq4baLeW7U9s3kLTQY5xL3XaeP55nYzCgjUEzYH5niDHdy3uJWY
KyHG+o31Nf4ZfTmVEzJLTCmsvvRpiSI0aPd/UiEHLV6syBTvwbmCNmPfPG3YGOFCVxkQf4jWMSONdcCnvfzvUCDTPDiR4tW6MjkiDXxTg6OUhLwS5X3SmID9tvSca+Jp
H7qsns+3drobOr+zOqQIWwIqMXIIVeK1r/QecCJRsJpObTw5Sy2iWiEo2KuFzUtNwsD2EqM4Z1P87X56AFCUgnWO6gc2PtlZPMa9D+dtFv2tCkeHPw9MIV1Kx8hmAk/I
rFvTQ7UNsu6xZXHZIDyxE12ZqFmu4Atfo615Vyf694JhJCiU/uxEu9UDk4UIFrYEE+xasZhMlW/FbFKVN4xzM7AtBEip6VSIMzNxJj9Au4QI5ORxFm38G5qLKIwfr+Iq
BoFh8IF5pJMfYlDAACV336L8rMamPpUrP3AmOY436sN9f0SzQghwx4RTLibu/4pGP4QUSSpbYBwYGkT6qqR8OBb2o9m6zJ0h8ltPadVQcPdB5q4tZV1hoaOYDFU40UVM
ENhV1iGHsuU7ClPkrTZnNDZhodOhr8OBOR3ZKL09GRO9HSDDV7tUMgay7EFEuhFIt2YfnFuJiNfBUOB9CHtei2kdcayNpSkkQs3ZD/b2fu/Mkc067bOnupePSV9zgwFN
MrTdOUwVnnkdRRvGKiEk4Z86c9J/S9a8sXxvOHzJOs38x6/FKn8G7XMx9HoZkzaLCV8mdQR7kpgaBvY8I++oGLcljhrIdVg2YaFJ03ZU/pBVLe84Ed5ks1rnGSSHRwjo
Pt+etkH3auOghj2W68uT13MGmRfno2SBNTVSQ4ZgZ+lrT2aLYrE8o94M8Rpyn9MAPh+EPFrh968odt6pDdRubsROmu8VUoN8L+0+wTm/tLai/KzGpj6VKz9wJjmON+rD
fX9Es0IIcMeEUy4m7v+KRgOZkBwsRQB6ONlu9q6JWg7zaw7UlHCsiFjTg//mId/YrFvTQ7UNsu6xZXHZIDyxEzKEirJ+/TSTR93gSFZrbLlhJCiU/uxEu9UDk4UIFrYE
vWgnmaeA19ADV6tfZMbx0bAtBEip6VSIMzNxJj9Au4Rxfyd2kRBwXklmVm7IeK2kameikCX3KeVwlF8Ce7ppBQzHywa80PrPdsVl+TBS7vAvcNOislCAvv2wC0lpnASc
wR7jFdqKJBTVFUu8ksJ9pyhSUJHn+ZLp3tctN1Fg5m9FA08H1GIFD0F4wfdnN22XFzV9LAjASyuZRGWWptkKv6GNDBt77KUCz/tuO4v8jM/JQUQsykwbjF3tzszqmmvS
DgRVfEw77Cs6TFHrm4htksIXIoiUf9ZZE+mmGk2bvQGWtxKnyIgQhjHDiIBz5H0bqpYTK5hNmd2Klzfb/6YEmYY/9cG99TuZtd+mJwW9I+nRHtwWsGfzGIhwCJGVBHgN
69IDkAoKpkT1o9yAMM/A7axb00O1DbLusWVx2SA8sRMH22Brn3oZlCQDW2EEkmxksmlqffmhtjRo1/vCxlhnnVxfbfGe77vCS0kuC+gvyrfOR4O9VmzFjVHqi8qqid+y
tmksJ8iJzVTC2bWsmMWun8LvWkCxRmn2lQYLixSGpec8vqlR1G62BfQpei9A6qtlLydfLPEzey50Sj2Zj/Y7P7ROYSaI8tcVGYdjfjOvYaeOSdGTPkCFARUEBxU5KpXU
4m6yjGtaNL8441cFffL3Nqg141JgOrHPLTp0kpLSzlJjHUC0nM4o3bKLJ46avyUgqIEkOH26tSb3deh80LsNUHik+ghcoRhLET/8nFyuQVLoXDeCR7Js9RpFSBqbPmCs
BOoAwkafqfZBs+QUeEgxlsP9khlfodYSYLBo4nDeULR5ess4VS5XF7cYqIZAdIfzonm2ClYtkTkXRqbJiC1HYG8ps54CzFuooI5/gjM53nOwzEJCiW7skGBU5rBPqs+U
/fBnZ5a31hh4nXdf4SNfAp8FmiTCF90lCl9I+aAv4YFRhzxZEd2g+oHxGORoAt/wyDbQhlVsr4GWGYK+bY/Zi7DuDShOS5iClsGrnQYwQVXosn9N2FkXyWaiqvpkV+KG
fVQXqd+FevgQ1G+y+sLtQnLIA+NbVZaB3KRO/qhji5tfzX/by2uc92z8+eamPaR8AcTvF8gwooMKmKArv5m08IGMHoZEMz+0hqBKnLDqUGfhFXmAbR6Le3mBWzt5QYgB
gzcCqEc4Ez0rMBh8j8egxJoFbwkoCBVsYFtG3NaP2Neho7kR3OxALiPCEkkprpMDlMfzs1cqN1mAtJ1jJCbSCIef37E/tspHcfFxESegejSonXee8WmwJLfVstU4TO6c
4SC6RuZnJQUeyc1PfMIVZhRohEeLkrWPSRsNwhsVCRYiueEr5TMpMFgWZLCIgE1DEuN5ItMR2CbZI+Uom/mcO6kpV+KG7ebJQBIkvZzjhuF0m4EEG9mVJ17dWE5OAOZ/
vRgkVrrMKm5klDNO3AbIXcu92gBjI9n4g7+WT5NbZP5rjkBAT4K9Fu0Qt/XM+emibN5MDR+1xUR6A6y9Y3m8nOu9iSp6hfStMsJxhHyV3tXD9a2dT6c49YI8/Cozi54a
Ioy3pLY04iaM4ShCw7ecCdLf3A8DFMCQocflX8E36B+fsYnMDb88t5mVwZIcDMv76SvJYmB7+UBBYGdUz4hNm2uOQEBPgr0W7RC39cz56aLpi1gpai89+h2BprA/kgr1
qVu6MnaBCMysuW8+bF32tMP1rZ1Ppzj1gjz8KjOLnhqQmuiKb7K3YnFtB4Yi+UB2b2c/FhwgFm76cayrLhJAP+yoyXdbjFRZ3eUZhlDfumxKwcAM3CLDQFtnnbEt0G2e
y53o8tnIq/ATSEG8jdEP1dNn9GKAMR2HpIqF3KtN3z9Ppn9l5Aw4aC52FIsRpNYKMtkqkbzzQ+PdBonCeMYcderfSpepYV7pkiMqxiIm7gVShpIHg/AIpZ7VhUJ7hkw3
BOu/Rvltd/hdf07jmjVfiqL+8sBAYnDeYAF5dFVjshI5s8kSv8aaJpf3MxyxvhmJjNrpVyXsPHTagFxhxNickd6m5ajH4eSjLc5EzGake0c7dIZlyj+GP8XsehcqYslX
b2c/FhwgFm76cayrLhJAP/yLubEocczZUw7s8UDiB3xQ4UnBkDIrATBm7se0jqV8bslXvNNJz15fR+A0PYX3g2F1d+3StbN3AmzTXDOcq2lShpIHg/AIpZ7VhUJ7hkw3
12jljkS5j4yrdHB5zYA1RYW+zQVDCQI+Vp5L1FXFLj1so1g0L3TE98NP4Wsr65ZjdJuBBBvZlSde3VhOTgDmf7JyTZTxAWplTPvR7xcfYOyb2BNh55TQk+b8gwIF7NFp
jZbR7cX1Ev7OdaiPXkm2hFpy1xEjbXKXRYx9hISkOKStlj5d1KQfiVjqiZJJY1NXpa5HyMIejsUxdC/dBq2aAcGvBlkBtOLCzXs2YqP3y76HfzqWJA8n3N0ZOskEtv8N
9pJOuPWP1SN3NxveOw+WQnJSb+CYKIJQEQgASFS3Z3I5a39oVwlTdcxCW7tiDXVM/DzrUg1uYipNlmUetozOg+j7sTTMtTtR7BJvXIASs31YMn5zIFKlu8KVM7ogQh3l
jH69aZXEtRWelqdfHpcjq8cpL0DXHViL6G800mKVJ2fTERIO12COYKabGTFtZBCxO9nLLMzYG5AmnOyUOV+VUzlrf2hXCVN1zEJbu2INdUz8POtSDW5iKk2WZR62jM6D
5xudeayE1OrX2RoXyBnbRFtJo5YnEfPuxj2n/2FrQjAzgKqy0483kALtTloQtRD2gP5xFWeckiJMADRAW20N+yp0RZtJIC/SjHJqejkldSJ78PjIYfo1Py8RU7HKBEHL
pa2i3OugnfSsXvkKYq1LHBgOYcC79oHu67iC+FDalVH2wseDjlzKlixflMncoFmdPMv/gKNdlvf/8Xiz/a/9vkEgq/y8BH5NAgW+B0S9vouQ6UtVgW7M14bMvXUewYqk
4KCgj9VlP0IWjB8RIQR8AQ6cTl1Yi1T7krHmRpuRMXz0GufBmAihKqX1pKF23ExCuaxmOrnKs+aDWQ25IaprxmZ1Wwr0xFXu7bqieK+8xRWiEkWW6+NxV8pwmZNRDnLR
AqWGRCHDeu9pLZlU14gqyF778Dk3CgQCFFRTdNLto0lM3VtS9paD5Gh0JOnP6rJ8zrdf9mRQYMPE5G13bsqd0b/j0zLsWmcgGGJXfhJPXhQ5Rl/2GlArZ264H9YW5h3q
PqT8zvhQq+N1CCyITz+B9Aq8hSniIs4tXfsS6diQiGZyUqNa3y+hg93v1c5luYoXH1pOwYXogUa9HaenTQG/5FGF+5bGyEQcHdHWYF5WU43cWtceiMRi7h9q3ChzO3+4
YJVNsl14VV3bXi12BMv2T+Xxhs05tOSe7UV1pfOji09ZehznO22FUeZQMBEcGtvdS6HEvrzzoFZRcksY45XeABiNc+VKLBs37vs+YbXaE5vXUvxfXVKE7CscwOul4jSo
G7f8jUCFH2gRmUjuHI7xC9xQ21gC7XIPfsYxpfyA07aYjV8OLeSUAptDpONnfU3I573T3Xi+NR53Jag+FDgxG424PkHsdGCPIHqVV+4+4fRwO1hbbWDVREueQDInwxTZ
8Ku+BqLjnoPGzVAlVCNy+EskhE9pS8LAYEtbY28Rrt8l0UBt1bMqKia3Z+3ifbRKYulIf+JmaWedyuMU9xZY8hJtYtFZVeWXBCECqCMnqEB5ess4VS5XF7cYqIZAdIfz
PT2qYPw6/mmnlF/3GlHo+wTHCo7w7xO8yp6zjPMT2xxW265UNEmEQPb7qKMprZP1W0zY4YaAPQWUTs1TWEQUn//BkVvHrHYYzvCxn0uAMdWkBR6MrbqsieYWviDOinCL
fcE64cehb+YlHsDauNvpPBabFs4bDKIECARLB75gtryuZh8XpnVO3HoJc7MsDVSlA4CSxgyMSfHZKbHQnSGqb1c0OGhGkwj0dgTNPHQhMMZbTNjhhoA9BZROzVNYRBSf
bD3Lceb+zjaP+hpw1Wv/naAUdgVhDyi0Wno0G1SF5fZbGXUALXTyia5idSbav9fvZvDPrs9hwJaMGjFso3EfY6kPFxA6V1E1e97Ec4bVkyIU4Pce9Ua+Vml3vHurfRvA
yogm0Sa9h4GMq195YwJtiHfjgJdSuLiEnmOI8obJNQoD2et9Th55Pmrxfj4iOFJejjBQ75PEGCAZy4xAQPPuZxThOEQKZ9IXJ7ZAGgEcrbEU4ThECmfSFye2QBoBHK2x
/jc8SLeMa5gWtxNTA/wsZdmdZ3Gd/iY20utOtjXTAVK/VQNZvLP/j4/G14neaAvVgvAefmJIGKqLYrycsKRw2LVk0uxyZzVtqpF6V8Qtu5ZXNDhoRpMI9HYEzTx0ITDG
Em1i0VlV5ZcEIQKoIyeoQJUoVoCc0FG5zuY9it+Z9pi/VQNZvLP/j4/G14neaAvVYiDTKAEXTkEpsvELGcccdtdjZlwkEumFTQKVPRiPUgBibuDieN6/6YLGJ2h3d8yS
lM9LFDk5XemfePQjdp0FiOsNq0FyB3YY6mzvSNNArjNIjvvsEbszX/GT89HSGzrEqjJqYyDySnealSXY4HKV/r0jlsyNsePw1MunTAze6BDSpvMHpsIJ7P7RpyH7EGpg
dHhWalG201yHmCBg6aUXdlcF6g8zfxKUcQ5oePF2bzflR0YrSpFMKwGhZzjN/KfmnRu+6k9KS/9uQT10PQ6gcs5oR2I2K1iyzuRB6WT0RF7Qlc64B+MFU9pxbl0XRnQw
1EZmFD40ajXoRQDlIbzO5mrB/tZlkRRN8GuVHuRFZCnINtCGVWyvgZYZgr5tj9mLIlaVhMopB7Qnufdjopi7Jlc0OGhGkwj0dgTNPHQhMMaqdGL1HznBQ640y/jnl+Pq
cwhC5Pk3BPO1DyVg0PB6zkjA4dIXmoXat/XzHmBcDrL2nYuNOcjZwYsikYWodOh/UeDuGc2ZpR9Qysyw9oIoohZLiLs2xaIcu6ML//XXTdhc87IOTcgLSaToZt+lYHjU
XGZQdVc3LCI2xQ4QvMYtETSwxsqfqa6sBvdlEJJOXvffeAfHU7Ip/yViPeljqEJe9xcOJerHEjE9H/SuWk5JtCMPJeykN9Ekrp/s1Ne5EnF6tox6npPn6JB41lj0ozK7
LGkW1xIh+Sq25ktZhNzdDJDqmZafgw82axBDkXHlkZnISqJTZmjF4hI+cxAs3Q+9ZI2+6MJGwutF71SRzls8lO23BSN9LmZ/pd1K56RKq7MptXAW/uWYgTjzc3GMR5LR
XO7hHnk/duC2aVOtdfWehgjqwUCOPDiGf3TKKwjhwVmb2BNh55TQk+b8gwIF7NFppYHf57NXehryHozM8LUjns/aggrh7aUiPQOdDO45dp0e8TAkIeHvsJg2vu/BwVsC
NA10o+a+EphK6yNEOLi+Z5vYE2HnlNCT5vyDAgXs0Wnp970xIkM8CExTRqTEeRQ5/vFC/UWPyly37eH05TCPiczuprQro/GSYx/SkVsxfKVDFeRIzeBtgo40QnRM20Tn
7PlUtjnAK0+gojtHjhfuXhRiwHZJEJ1ypqqKgExMB/bOkrEF7cMjb0Y6/INvWCf+kSlfj0I/haoFEuyQABotJN4I8ubpKt7IJYSwUTeG3Lzcgveeq4JozZfpz3rzG/C3
lX33y4cj1f99eBOMW6a0ksf1uwELhkQNJCv2V7wO3Z3K77RB6IEtqVOQ2ENBHstxV0qtsc0oR7X06bTRgur/mcg3qYWSDTS96GAsTXxSfVoe8TAkIeHvsJg2vu/BwVsC
Q67sp2xfE819MZJSdI+XD1gF9GkqvI3T532KH4N1qB1+FLqUoYWgfB7tzHlVe3fxREceZrDM+j15c42TnRvDTTs+FcowHIPWZY/nMBcBQ158uJpTqjaDMZLsDmEKTsFS
lmTBv/Jsyh2wrXC7dMiOos3OqvbosFkAM/spQ1QrRbIGmx1Wdi0ifX3CLrdAnM7ypXKHsJV0YqrkbXM/od8iOlasp45qsW82X3LhYk5xYCgH39EmOMVMnxKb/oAbdJxx
62sdUJBGmnwIAri7z3dXY51O8B3WZneSzlZYHdc5WZlkjb7owkbC60XvVJHOWzyUVeXeDswjPaUSpJtBLm7MIkvBIBLse9AOzVQbP0+Ib8yLJ2V2PvCiEGEO+KqrUptQ
Jbci07E+Ls1eMiqTXYNG4/ifYfiqLxgTAmEGvzI+TvfZg0vMoIo+NS2N9x+CFjtzyLVZQN/7EUHvj2i78gkCc8bqxvpb66XJKdKn8TQEjC24r9HCeeA/FAShgYiy6oNv
qxv9SopsaJSceDAfPRCdl6NDS1xZS3zodMznQ+6mgxiamVEDrDvaXlXSjfiplOZwMxvYJpvEFmVIuQfTwi43losnZXY+8KIQYQ74qqtSm1D0DS0sb3hTKuz5jdXshMWG
3vc9aqxMGeFpaENZyuJ9gJO1h6rFMizJ++C2wMUhGuJcQ0P/+qQc9Zll0CUSnhLytGod240Fg0uv+Obc5Xqew/W3MFAzdWZ2C6EXeFns5MZYBfRpKryN0+d9ih+Ddagd
r0QmjCn2/KtuskejV8wFH8PjDqyHPx6zskyBy0Ub3OegXZasQWUPvZMsR/cf1fCs6l892WloiAwbAAPeOPKzcFqEQLSwtsnCpxLsBBuidn/eVNoyZzJgIwpx9HhbqCT/
HG6P5l6MmxnGs4pm7iPzeC59ndjpPcaMq6uCoZUgT9LrNc2aPiGyL3tSMALfWnVw6u7YhKEvUT+clqnkL5IMOaNDS1xZS3zodMznQ+6mgxgMbzAjFkOMknarnpVRO0do
2xDCzfjQZp4kwAcvN9bD9RxxZi8K+Hh4vJxjWhSX1xPXNrVpHkyYZqCvfT8EZQ3AtvVpGoJWHnRYEPOGUh6p5Ylgk1hC9b/ChFEkRsxYp4tYBfRpKryN0+d9ih+Ddagd
r0QmjCn2/KtuskejV8wFH7knhvtI3e0Ov8bzKPC6whBtRkRQykKm6gTvzKvgUS3kgr+ZygLZSJq8LdnJKVDHsb4kbrPNdmJ+3mjeUC1JXzGQl7R1G73J1Kx0A556GbKO
qNIDer5oANwjitzGdMFNTtkUkRhUpu1xxYYmXZZgJO1GMiEI7UqKuJiVZUczJAOIU5sfrIsuBQu+vYP36m19UN2frUoTqVGuLRCppXr8f7yjtOMI9wF2UYlJYrxhrqqT
IlWJnguEovWVZNztjgwbrxOMZefDyVApuH3NlGV2gyfpDwEEZvyPjqh4KSNVbSCovpP4kO1fx6PUz0G/FZb9XNCvExSv+QYXYXcNmr0atPc5Cf7PbuxpOx/n+8EYnKzG
GwlwGoANGGX1DlTUA7x7vr4kbrPNdmJ+3mjeUC1JXzGQl7R1G73J1Kx0A556GbKOh63IXSrZoPLvKd5ba58qf2SNvujCRsLrRe9Ukc5bPJTJQFgznB3khbuGz0lAm0ac
yLVZQN/7EUHvj2i78gkCcwYdTyCH4mR1vvygUtKipZkVPlbhlaSW1dBikFqh1HKXxJgT0pNCgmeSk1QS4wGXgTyc1hfKpU9moQV/he8h1bO7DIXWP1pfviKyhDvg3Hxu
xurG+lvrpckp0qfxNASMLcKDC0hqo77A93tKbBovUeIQiSzkvh5Gw/r3o4FAFGHBoMCTDUeHrEU7FM3Ln3Y8Cwin5zd2t2uGAPQbEKcYilPCuFEl690/B3jzSHMHm4NB
JSVm+kCtEEXyQK49qS3KWumEkVno/l3yPuzG+t96/Na+k/iQ7V/Ho9TPQb8Vlv1cIfLOYXsFliYB3Ig1dSr+/6iUZUq0r/px5W+qQYIyYFWwxmK5PerJY78bP1LBjhZx
xLl9Viujq5ehDnlK/3oa4hxZ0c9jEHXy4ySPUSaCHYVknubqUzHQ2Cbcz3aTJjg+xJgT0pNCgmeSk1QS4wGXgTyc1hfKpU9moQV/he8h1bOC/fC4NWqsPAFMrnF4SFWY
SNCQbyV7/HV4p8jjgZdtfnESVqJRmzOmOtFocOemNatQ4UnBkDIrATBm7se0jqV8HE6t1dTGrSYngr6zsHvZiwe/3n4m6BaRzXXDRVYafpBrjkBAT4K9Fu0Qt/XM+emi
iTGWiPds2HbTQ+oqXmIbz8BHGkdCpBEVFc+Y9V217TzhJ/GtpzphEEFLy7/0nBZ9iLtjZF0L9QcZsyRvbALWvstNAprDKFZOrSrNBnXaZRujWn5NszG6EYuDv7tyPoVk
57f7XTgsxZ+4rFULRReop5CXtHUbvcnUrHQDnnoZso7KqD8xF2ZOOlnI273onR1COz4VyjAcg9Zlj+cwFwFDXoVTLGkI/xvhNEulUeuA5t+WZMG/8mzKHbCtcLt0yI6i
zc6q9uiwWQAz+ylDVCtFsgh+wWOIfbqgTVbHOfXcLFGS66GGriZVbWQMaHq1QE3HhEU91Mpo58cS+nAtkLDJTn0TtHxwqJJ6OEwPjktvxqe8eMDU3kwq8F6AsCz++QZz
TguL8fR6CYOigAGnV9oR0MrgbPwUUxJelkgpAA4ZDNM5Cf7PbuxpOx/n+8EYnKzGKZWiY5Yb59HOzWLtsjojNkogazM7L0oI5486ec+sUNGLJ2V2PvCiEGEO+KqrUptQ
dXiiFyIXXvnxXwRdYNgAC3PzkoY4J2AwZxy4yEkdqpEyPV0MzaFVzmY0yq+rD22cxGb8kLyG5sPxYcyB2FUtLVLHolebDXbIldxnP5shBNX3IhSO91pyc+jKKzsb4zxq
c/OShjgnYDBnHLjISR2qkYF+GUsnBAH8lKneVB/P/l3oIJdQz9nzaONcUARhyhm85Fc5uvP7rDNROSjdT1Kyv09YB0iPByVrbL05v0Q3uiQQiSzkvh5Gw/r3o4FAFGHB
fhS6lKGFoHwe7cx5VXt38Up4LaVSXiFPwZeVoTLQfUihDV5ehn/+lVqTOCeMfoVDt3Xo0A5gGNGA5T4FFGRJDfDDwOLm1IBlmRRm2RwKTTrSC77SyJmCm6nUDYygl8Fl
b45DJQywtyOzL1VoDZe8X3Ma8hHKM8TUi4Ut2A6RVjaHBLK0fm8U959WYFvepcBi4XvaWSRBvIyz7fGBXo8aeVLHolebDXbIldxnP5shBNXFVIBN4MSVMhUcOR7NT10+
xJgT0pNCgmeSk1QS4wGXgfgwzH92yJ1yY96Zs7RW7QRS9lpp9/FSoLirTWbertxkHQ87wozU++4tjaY5ADzpvOD0OtRV0JHFkkWJNfnYVqEQiSzkvh5Gw/r3o4FAFGHB
I6hXTUvv6KBrCduTj7NNhgvvVecoDsl0oORmQgFEiEdgrL3bOrjUJ91cgceBjQiLJS9kqNFqwWOXQOIy8LEFg89YWInS4C5SzEaHVNuYCSIgafMhFhuHbn2i+Reiu1ms
2J9unDA1YdSFgeiW+PKKcB7bMSAVSILOJZswQ3IGStnrkHRXQf7FAQPWO2Rp81l/m9gTYeeU0JPm/IMCBezRaRxOrdXUxq0mJ4K+s7B72YtTzY6GKOscg3VBZM2TgUB/
HQ87wozU++4tjaY5ADzpvM+oWDsWGZERYMia3EhsRToNoLFGfnLasQcS/2kzJmqLtrfXr0S0iPm6dmTRE9m5LlVzJibHV2IWp1FasxywdxgdDzvCjNT77i2NpjkAPOm8
rxckGLhLTTp91WYCExKPqGSNvujCRsLrRe9Ukc5bPJTl/nhwjT/CZxHFlV6LRSr2klrXCU8lnkJ3z2Y3tw9IVyOoV01L7+igawnbk4+zTYbA1q/JpR3msQblhXy49od/
xqpDgFqymu6ZCFhJ/bIRInyHPixWIgAWOGUBec/OeZh+EOwH6ht899Sijb63DRiqyLA74Iw2FjQPMPleeJ4vclEN0XFVS7qPH/APwydBTrE/gl8dff9ijRnwZWzNzW1/
fLa7BsW1A+XQPlLSMlhNj30cAOAiKMCG7wkz5u0MqFggafMhFhuHbn2i+Reiu1msr9QsWLdQuzsj6jpaNSqQtT+rl30tmBgXrwVCsnyrrCFC2SZ8RS0ftOftsC5mfZf7
p8hWchgU7Vem+xDMWw16FjCiPdZS8S4wRBjkAWbYMRdFY2iEBMClLkiZygefXHGNM86kYKw4D6YeTkOfKOwcsn5Zh4L9P17P/Ue4R059z8evmrRfp3nrzYDiMWazyjn7
adQHe9rZNvBVfeNlmdsWniGhgvOwEoAcODwYWM0UC/EYU02Nae2KQhErGW6iA/AJpgeI0frX4Of1tvxaB6Fmkyt4yzJRwMwbtPp+vPYF5BH09CNu0+jjp2LNK0R5D1wV
GUnjBL5htQABe/EhEMqv8YVzV7gsHbzy793rofuyKxHSC77SyJmCm6nUDYygl8FlOe5aBU4e4w+8OGLY3gm7Wbf6lUuLqv9w3k75tL26zwPvankBLcwM/i9EY/r2Oghz
HHFmLwr4eHi8nGNaFJfXEwxgPFjJpEG/afkuVi56AgGAE6mQlh5Y17JyHnhl8NcKCgy0NKkAjaL1LnsSPycgefT0I27T6OOnYs0rRHkPXBUZSeMEvmG1AAF78SEQyq/x
tnXBNKwgJR5Or7Za8ptR1Bai+qM3N/BWtfH8tr8WTPev1CxYt1C7OyPqOlo1KpC1FeS+9jZPWWn+zZBJLQH9JF5sn6XPeBngnrXCgyJf0+mo557DH3MQ3EvDJl8utriu
c1Wq2SfQ/IdcTX/XD1fH0UPdzPBj7MY/c6uxffQEM802XUTZy4bNU61F8UL+rLiBNxqE3oOYkdgHDG+EUqBkbAhXKTQ6nk964bzz7PxYwfHCeGlVO/DCgmv9+0YTEOIT
V1EYgLhHB4eMSqcK90tPmmJzCKKWki33tt6f2wDIkO+Q3U9q3FAufoBEPwYYR/v1J32dfO0r7KTmYgsAKMX33rRPitmyAq516sxogUIJLFheEZ/uaKQpV5/S16Wur+ba
FTElagaODzA76YH5+FUtJ0lXQ+GRYKordTkDtdaestDS+NfiEyCHjJj/tdIYhOYd5o2GRkz6ceXx5Ax9dmnkxokX9yolj8/6R1j7soxeXk+X9/SnEbS0v3WJ84P0/ffw
gkLYrwD43wGbCfZ9vwDppc72vEozHW7KMEsGpDYp6vpJV0PhkWCqK3U5A7XWnrLQQAoFQrVutPLQ+As0hQn/gMqIJtEmvYeBjKtfeWMCbYiJF/cqJY/P+kdY+7KMXl5P
r5q0X6d5682A4jFms8o5+9t4mowQsID/3OY/vgLUyGsxm2maL6GlpYiRgU5p1fFlPU2FIchIHgDRFUpIu0hFh6yjNiyQ32jyO60OL/DyFgH4sABhnZKlgB3P/uuyBEIw
Joo+TJu7FGWrInsE3nUHJTy5wUiHGMRSBTDqketQ00Ktlj5d1KQfiVjqiZJJY1NXC52cWJSerqdzx5thGAwVNhy2ix4FwUzbMyaPn9APi9JPDA7oub98bVjvgG+0+nMP
U89LEFx9zFW7Vd3Gc9B5SkvvQFVaO6TIL1fp96qVqc4K41IaCDDFXJQ+j1FRAEcr4Sfxrac6YRBBS8u/9JwWfSmXo0c42TSUYiORmpi7lzLjKXvm4XLKCjZG8NhSRGba
sM+sLOC3yGjoxPGgBo+9id4I8ubpKt7IJYSwUTeG3LyZF3EG1TvYOsmSsQGULznqp00ba0jt/DEiK5K2Ee6xL+trHVCQRpp8CAK4u893V2OYwMQnkHbfgVgNlXAg6A0Q
IVKyrxFMoqVRgAqdJCjFmkg75Ye0HKEzWEmbB55VD3YWAOWCELPqYw3s9eqzjt7lYiuyGtT0ZojIe84PomMMdwX2hq6vfxH5D7xk7LHUGWcdDnDV4VvQlhOsqttR41jm
Qk0iQGDy3UQ7RCG6A6N36hlJ4wS+YbUAAXvxIRDKr/E+T7BVmK3L1gdwB36mEpToRgm8T5j4ftI3YK3axnR+UyziXmBvknAqDzwqJMKGTuklQIQUfhNc9A39rHziSDru
C6A5qpX4zaD9YzP3omMO0hxxZi8K+Hh4vJxjWhSX1xMtqo+Qha/3XEesVdITDYhftAKtZfxABvorZhN3YIozxyc9TI8VVfxwqk77JJv5rch6GpT9GyK94Kh7jN8DadkF
fLa7BsW1A+XQPlLSMlhNj6tFTXRdsCoVPYAfaPW10HFrvmfC0bStZKXmrVGhpYpYLOJeYG+ScCoPPCokwoZO6RwSRd6Om6AA83OJ7vbVIl+bPHvIjiIERCJI1GH5BP57
3gjy5ukq3sglhLBRN4bcvJkXcQbVO9g6yZKxAZQvOepa6aUKufAb0zzGn4rntwbo+LAAYZ2SpYAdz/7rsgRCME4vB/GvDvB8MEHfKi5rRtiPsK/wN45TbsVINR5bLNxi
MrCduRkzylrLuSoMOcjgp364dE/yyJh/sYkPUmdLvBWW9l4QIzGATebv3zq7OdS0Q93M8GPsxj9zq7F99AQzzc3OqvbosFkAM/spQ1QrRbLa/7amaBLbDIE1iKuv+ATn
2vbdjv2ioZ98CAOGZss4wp5haPN3PCGs0MVjW3HenbzHbgUrs/bvBf8vb3uyI7LLyLA74Iw2FjQPMPleeJ4vclEN0XFVS7qPH/APwydBTrHQZEMeQg5Ld+popDx/WuW5
FRe8MsfaJ/3lhUEcM6pUCYN/qRvhWwjvKE0755rKsOuvRCaMKfb8q26yR6NXzAUf1PpYLITXrgecYUhsk66WvyJzZXopwKz2ddQvTTSeVMpHbE8R0jHvFGkRAPbPyPGB
gUFKnTqDdDIV8b1OjXFxNhlJ4wS+YbUAAXvxIRDKr/FnPDxKguON2AecB7LhOZM5Nl1E2cuGzVOtRfFC/qy4gdr/tqZoEtsMgTWIq6/4BOeOSx+f29jI8vnF/dSnWDGD
PTb4bmBcd5lMtSNG36CzfAJ+VBQL50o4Jq9FdKDFLFOCx9MdnR6irY0c8+ETT+obDyTFZE+koBq1JVGxGMCzP+P8WLQHPFHDjnRKnNPNsxwr7qZX6//ardjeGERThQkG
6+2BhyKwcO/WVVzDH3PYzyOoV01L7+igawnbk4+zTYYdOZ91hJtopV54xeH3pHnfaPx7CCqD12UlA/I89e/F1mu+Z8LRtK1kpeatUaGlilh30KAV/l+/57qTi7WaQagi
P6uXfS2YGBevBUKyfKusIShUcgoxtL5qmxVnrMJ7+6bg3+b0HEdDXn19kRpjKfKcGUnjBL5htQABe/EhEMqv8bmacS3wfo48jStfhoSLIvs2XUTZy4bNU61F8UL+rLiB
d9CgFf5fv+e6k4u1mkGoIo5LH5/b2Mjy+cX91KdYMYM9NvhuYFx3mUy1I0bfoLN857oRgMZBce4RQWtol5mCoYLH0x2dHqKtjRzz4RNP6htn5lG+bIvb/3t0PGiF0WEb
qr9G3lX8tkxqBqg077w7ktCy7yKV9rOVBTDcx7XEwrTZLLGiyuxqyjDJRhKHgFPHtnLrvRH2pLTHIoE9X+pwzpH3X8R0vLpx4zYsztI33hHKiCbRJr2HgYyrX3ljAm2I
nkPELMSQBI3KYVRngPExRmg4IUyvv7eflm57V36/07oy4cZoWKoLRVrjQc52GLJLNxZvd5XJGAVMmoQB68QqHjJI+fmFlG6Fl0bUF3LVAo9PQB1KjT4ijF3ek5qmB5wx
UAwbLiqqh0viIfFExnoOClnOmRy3it6ooBLZt9FuVpa4YWjxaqk39rqDGQqHunr9EeC7kPmsKMQZKsAumoli98qIJtEmvYeBjKtfeWMCbYhQVwys3bC5W1JiegIIlSi8
5+m1y34Cg1oZVSyTECKRuQvag6/RCE2tfJOzVOa3btAw/QtFdEmQOQm1dfsPf7N9yogm0Sa9h4GMq195YwJtiKBTe4B3k/mbHjIUfqo67SLONWsHuDzSUPpB31bSUBQ9
/4rNcVs/JXWe0ojiEfKz0kZaWtRXrNKJKuYfu2c7SQ4IHI89GHO7Fgaiqszij2Yw0yGRnPZE1s62DA8g752IHL7Mbe8/j+Ht4dB91ap/2NpfofKWQIXEJP2gAPwXUZ+p
KtHHUmYJBzO9SUDZlVA8xElvLRIDcIs4P2iBz5rE8LnKiCbRJr2HgYyrX3ljAm2Id+FUBXZ3L3OKxqh0id+YDJ0f+iTMWSTw+NfqdGf4OnPVbSlwnefvItbi5hVpfOEP
C86jAyqIJ6dlVR3SJOurX8qIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOejCfNcbnQ8eC8VC3A/6mcJ8Qr6PA80SUB7r4NABpOzmUT1m+EkwmYrki/Sk7jdQ0ov
Y4so381Uz16xW2ffSPriyXIHLql8/FShcQ41SVHzY3afXgQys4k3WpaJOYPvlSAxAOABJeKTTQseOhyzRCxEw9CV6e7ZI0VvC6SeUIj+Ok9LZYbFM0g6MB7muLpZq2YS
yogm0Sa9h4GMq195YwJtiDpnAWVVHivKDTBw8yw4csFIWuzDG7iBv151iF8WJfeWa2vTfUyqyLiOj2/MT/3Ns6s+xqnRnNhgVbdMAbNnFgLKiCbRJr2HgYyrX3ljAm2I
KbAWmvuvd8ilV1icDV9dy8BLGX1UQGGlSBs0L/OYhgkkm8sG9vaymH2B0oLbOncLl1TgTWvMurZ3y1ihSz5NdG49yqOPgox/MoPbrhsZmZ2DcRdOfnzDCIY08vsxLu17
lKkOv1tpoGkegjZpOahEEBMjnGxcF7FoD4asjxrz2Hq4YLHcDzqEbIctirmY3/dboB1H7eess8hzaBA0sl1vHMqIJtEmvYeBjKtfeWMCbYg6Cy0VxXZenqBxkRlLe29K
pLxw/MtCGNc+PS9CUXgpMvUOzgVhr2GoovWyiZv7yBxL70BVWjukyC9X6feqlanO3fdyYNKT1Io2V6H63wgKoUDJqrCQCDOrgCkmTBNGpAyB2W64YNcn0a/5LnMyYUfj
2ztesKxOGtpVarBZXHKvN0A1vx2RcBKx5BcgBNPUegzKiCbRJr2HgYyrX3ljAm2I9eAhsbYpcvuVPp86ImPIqlisWByskj5/vDXqZLmdpn80zmEreZem7mOSLCVFaxjH
0ydpNqWT2Kv1z3nbA/+rMhlJ4wS+YbUAAXvxIRDKr/G08H35oy6GwItvHhk8YumWaE7tq/7wib4HT2wPH0lGOLHjOwuJurIhc/irSU3VqEm4UX57pNWuygLzbJtmqX/w
LaqPkIWv91xHrFXSEw2IXw79tZajyFDom5bCP7KfyXKqXU0HtT+eMVTl9oJBjZfX9C9RalY+QmXcGeaheutH79xdrCTFVtfQ4zeRkTYrgKYs4l5gb5JwKg88KiTChk7p
NAPeXugFDkQS2Len/uXAB8iKr4olDSOK40NKSKJnm1zOME33e6e1TCr6rznNWp7LzigbGXFeuu7Hc7+UvANrPjcWb3eVyRgFTJqEAevEKh58trsGxbUD5dA+UtIyWE2P
l3rLg6o85yqXYD++AAzpQBdaBhN59OBztKdEqNin52lbcENxYwcIFB8hW8SCEFSUuGFo8WqpN/a6gxkKh7p6/UlXQ+GRYKordTkDtdaestArc9Mt9W91pmH/+SFFLcl7
pVd3zd04KWktD7F0hC+Rxu2I/CcVnwC/06ALY88iEiL/slq4fLX58qPt/DjN9NCzKZejRzjZNJRiI5GamLuXMne6iy91hKoNnehYFsPjr/mT/GB1DJsNpCJB+R8joIsv
qmvt+9RJG29CVijnCj5p6jXMVjSjyOZnXePUuYOLcytpO04tMhU/z4Reg2f08ucVFRe8MsfaJ/3lhUEcM6pUCenkmWUB/L4Hg5Kh0UN+xWbXXBAC6Vx2VUf6VLxt9KnJ
Au06ZOBDJvvzLrHj4wVs3irRx1JmCQczvUlA2ZVQPMSZF3EG1TvYOsmSsQGULznqDVLEMnuAhR7dW0v66M/gL8a1omAuN7tugAFrz+M154td0q4SXl5z3eJ5hapBQiZu
FOAnLeaNF/Ymkft7tZkWAJlzsW3iA3DBZj7qDDVptuU9MMPrdwpbidNNAAGPZlazw3/iBQxkhySfOon3kgYTR6yN31AZvu06PLFG+4zR/9THqzBB5Vi8q2TCc7/axwm+
Ti8H8a8O8HwwQd8qLmtG2ENoLPzK5UFMvHE4Vg1AzLCD1rGsUMNU4oi9/CgEJ+DvaxF6wE3QG1oGK2Z1Lp01z0RbntZbeVqMliJG2TRMHHx43JB1o6XvGQpgmksYx0SD
OYoPaBl8dJk6FZ6viaesm6+1iEFMvDUAIjdRH3DWCWGFHOcwFzwhTqXeXM7xhSIU/JKZw+xnj/AW5DS10NFid3ILjpckxD9y2j3EhJVZVgRiK7Ia1PRmiMh7zg+iYwx3
3oL1ghR3Pyf/u6aNj+4iNImvX5jRYBoyP+S0/fQvdRrWo+c895h9TkFlYZf40xs98O4WkVNhSDxFU3X0RGc3i8RsBSjK660L2SVpHbj0cSzKiCbRJr2HgYyrX3ljAm2I
g3EXTn58wwiGNPL7MS7te73eWELVj64gkPJAtiNhAfzP45sqZ4YalKRdnWUMnbqaV8jOS1muUv7ln2fc45H99ic/zDhU8lPwC5MfkEe7ZzrKiCbRJr2HgYyrX3ljAm2I
SjK63YNrrsokUjouvmThXXeV77s5eHXp+kZ/4L1cJNWlEGXn5EpV9CcofEFEDkTvCcBvhCSt5lzzPQLIGQ0EpsqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
bXpZ7ZFI3m9DByUulLv8uo7iQ7nBaKh+iDx0aaXgHgCAo79L2BhBoQd4X80WK8R1yogm0Sa9h4GMq195YwJtiJQcVJWN3VgEeoqzEzbIFtEiESg+1QgNvYVq4Dqvr5KA
WcnJVBEicAzEPrVJOAkwahBo2kHd8ilICKOw0cvac0DZLLGiyuxqyjDJRhKHgFPHtnLrvRH2pLTHIoE9X+pwzvOWPCsj8xBc+j0nBiPszafKiCbRJr2HgYyrX3ljAm2I
gRrInBgZD19HN9j5BZzno+F0tkNX5wrUi2d98E5QWohTDleMwBJM2464N1AuCW0vJoo+TJu7FGWrInsE3nUHJTax0AGZEijTPV6ZA2T3Kxg2ZZaDXYXXaWDgGk1XVTzH
ePZFTcL1YSTzMixXGb1x4P/iG5Hcq0DDyBJ720sziLHlHP8dyDpZs6MLbtplZyALvdDEE33/Y/o79/QXczL/adMhkZz2RNbOtgwPIO+diBy+zG3vP4/h7eHQfdWqf9ja
Yw6USLaMdetiVxRBYN9GlWX53FegRaXhBoQyRroTBzbI7SJF8dBkUnCj5bht6C1Eyogm0Sa9h4GMq195YwJtiDoLLRXFdl6eoHGRGUt7b0rjwzB0dESZMad+ALHT564w
ZxPT0Q7Z8AlZzyYu1Hv1ujBfPsc8MZl4v+tsorrTkBXKiCbRJr2HgYyrX3ljAm2IUFcMrN2wuVtSYnoCCJUovDZUdEifQ1myNbNn07Kl5YQPPV0IYcD1ooRMQFH+h/vL
9r21GyGuDPGCD7eWQSjt+8qIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13LTUWrZfw8PKnL17Wkucdyw69vykohQydzzoJNxuQu37O1GE0b6JLm4hSzDp96ruQU
oaEEGJs6RlgOQvlZzd69FKGOGRbTFlHiOvUQpjJMgs1Sgo9EwxalqN7NWcCGUv+52IxgPx4X0/eBdEw8eySRiHk3EupRC7Kztg7iIdy3O+PKiCbRJr2HgYyrX3ljAm2I
cgcuqXz8VKFxDjVJUfNjdh+Kt423vzRqWnLCfEq/t6zSdhbobVdBNF02DEO3Vu7YnqK7ksOLuvdd4fVhDs3UxDCiPdZS8S4wRBjkAWbYMReRFNRCU49O7sIS4/aqV1ko
aE7tq/7wib4HT2wPH0lGOLHjOwuJurIhc/irSU3VqEmfpdh9LxaP4kNirnI6ICLUSVdD4ZFgqit1OQO11p6y0CYS5IKbrlbJOI62qIqzT9vGtaJgLje7boABa8/jNeeL
JUaCo9bHheyTXzLc3/Xiv5XR040xbmpG3HZ8g22388FzZF/TeslayEN0KJnPX5IEctkxgQIXWav13RYykVd89IkLsgxlLDVhN/FrX1nIQ65VhXT8lqyExqEbA63tf6qG
0tL7ikQCYLhCWttVRcQn7efAfIvCERXvtTLZaT6qirb5T2Vl3FUH+2E6pXfW3xhb6cdV+3ONhDnp7Kb9AzvcQtigb6tB93qfUVDmIu2nn96NT1ZA6k/y/vJI5VlWNDkG
iRf3KiWPz/pHWPuyjF5eT4+wr/A3jlNuxUg1Hlss3GIHfc6gwaodS/rASaXSxs16asmkeyKg3f0mVbEndWHE5K9zhqSZXi+R00IONtoVZtEnylfclXCR+ACTr52AVhha
j78mX+Q9yitlyF6miv01E4u3Unb3CXRZhCZB0VExuKwG8tr6XNYiFN3irGxv5rA1BoMiHPw5GySYp51IAbs4wXTk1xHV0p6uQP5tLXFDMVDKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiM0IMHlIf7x/msBKJ2C747OAo79L2BhBoQd4X80WK8R12xKVbWglVvs/Qum5AlqAts/jmypnhhqUpF2dZQyduprKiCbRJr2HgYyrX3ljAm2I
0vZ/C5D4uxV8hGR06yAxc9yD779f3H8IKQ8+YcxHmQTkInEXnwPC4/4rNc3ldMDD8PE9HfeamS6wltAzhIgxUMqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOej
X/4kxAXy0+nESnWFF+Z7lm/Ld4unKZckBlhM627oUnXtejqRb9bd/j7itXgW90/xyogm0Sa9h4GMq195YwJtiJQcVJWN3VgEeoqzEzbIFtENVsRdyitV8jgrcL6s4KWr
a+gc4sVp0upA9u1KEVcZFcojENZqBMTUzAnLi1JP8ztUT/zAqMvCcW0m662ubCJA2ztesKxOGtpVarBZXHKvNx8eAvztaw6KWrxJzNedMdXKiCbRJr2HgYyrX3ljAm2I
oFN7gHeT+ZseMhR+qjrtIkBt0wzrEHKGfkbnTxSPWwXfVvMNN4aFZPRb6ILq+974CrS8LNpvTI6JLtBytxZJv5OoGuZA4Ihy2mJE7wibcmmDcRdOfnzDCIY08vsxLu17
nkRCJtwx2pDA8iXoCiLlKtJ2FuhtV0E0XTYMQ7dW7tgw5uVGUjzlaxPosnKc4z6/wkwFEbevcrsf6wFGLHGx4k9AHUqNPiKMXd6TmqYHnDF9NprB4chgHMmb1U5sOQsH
eqkudvE5PKF1wbyxin42x4gfO3BfgA381744N7i7Lb0DkGSLe8kPx8VxMZfCNN+Syogm0Sa9h4GMq195YwJtiDpnAWVVHivKDTBw8yw4csEcWwTuxn+8eHMLeIo7FyZs
FmwTRH5xaCll3M4ZYyNQqxjeYSm2VM34dabATX+7JjHKiCbRJr2HgYyrX3ljAm2I0vZ/C5D4uxV8hGR06yAxc1x1M5dlAwGW8ut9rog8Hve2cuu9EfaktMcigT1f6nDO
2v+2pmgS2wyBNYirr/gE56S8cPzLQhjXPj0vQlF4KTJ9SChKNknSZ8s69N+tqhXOgnOzlbhy1j959VH45Izi9FMOV4zAEkzbjrg3UC4JbS+Dc9e3quubzCHoEi7ACxnq
yogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKpYrFgcrJI+f7w16mS5naZ/hQO32xnESp/xDrB+UEDYYPgu6vfhrulk6OSvvLkEaxl8trsGxbUD5dA+UtIyWE2P
0PYmguvD1iR3rNo2RU2TvddcEALpXHZVR/pUvG30qclUNnJyF9rV23ZSA1cJGDeYpivL25oh6tmzPxN8N2x+nfME4ODJz2DUc8v7Gusn6CdXC7gsWVVP6wPjihBxYEsM
6HcqaiYxO3xdTuvKeUVmXrIGU7AMP8ivqQkYl+xtL6H1Ds4FYa9hqKL1somb+8gcLaqPkIWv91xHrFXSEw2IX+vZnXZy9p696bIWB1qAsYKlV3fN3TgpaS0PsXSEL5HG
SCKAg+Qr9pGztsmcjjHj2GCrVZDVqX/iwSS9ZKr0loa+DtkFneJ0DY3DpZR1YZcK9cOT3nPi68WQpVuOiiHiFImvX5jRYBoyP+S0/fQvdRq8wNfhDXge6wiK0QpZwdwg
6s/QiXqzNYZYuh9z07m7CjmFbImrX7fv99Ql3nZjDcgu67PhQQIk+j726hBlMYDGdHLXggq+2jbSssGOE+nMeXTk0Y1LUQnYNG3nEWRPfNMJwG+EJK3mXPM9AsgZDQSm
+VdsQrH0fz5O19+O491ZocqIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N2ZVkpmTsX3TZxWewP8EXy67P1QS+NChp/5RRIpqB27DBHIFSHfejkKTDJBMTEA0sa
vkYLX/miMK4iRpo4KSekV94ER6ENG7m0FDD1bgBFTDqKE7BF83oZcma+AUoggFGolfp8vto2C4AjUU+M8T9/EzgocIa7zk9fi7SExy337OWIk82ngUM3c9mxfKXeXDQy
yogm0Sa9h4GMq195YwJtiJHy8a+t65Pgk9YYq0n4lq3+6KXMO1XMb+/bBh0zRJ0FQNuG1YF0DMQaoPi6gbKncjDNFD8gQC7qU++CVTMinizKiCbRJr2HgYyrX3ljAm2I
q5EJeO5pbNbXGZg7gN6EfAVeEVjpIyRnsbM+CLRSuoGIHKDIGPxpJBl8zpSWasr2r+E64KATNK6JX5whNyUrKe5Sm4fRDe5cHPex6N+Y8I4opYIO1NLAv81sj1hVgi//
2nwprEjEJ/BEkk9longSKcqIJtEmvYeBjKtfeWMCbYhQVwys3bC5W1JiegIIlSi8NrHQAZkSKNM9XpkDZPcrGGCrVZDVqX/iwSS9ZKr0loav1CxYt1C7OyPqOlo1KpC1
4/j5DGYCmQ5r0e3HF1EWw+nHVftzjYQ56eym/QM73ELONWsHuDzSUPpB31bSUBQ96veHphH2GpjPYNYrlftWAO/+//3zFuBc6hpPyFOP3hyWYnCpLHNzGAC4XS62ftEe
0yGRnPZE1s62DA8g752IHL7Mbe8/j+Ht4dB91ap/2NpjDpRItox162JXFEFg30aV6LHUMREqEBXOZLt6guyLE5bwzClTy4XZndapCNNU+PPKiCbRJr2HgYyrX3ljAm2I
d+FUBXZ3L3OKxqh0id+YDNkZl2P/4hmU5Ym8r/Hz2EJuJDcQJlFnPpeoikxCl01Pt0w3BgnPdKpADgobuDZ+ocqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOej
CfNcbnQ8eC8VC3A/6mcJ8RuHtOR91HElpuFqZfzwZibRv5n4W+QwCGZG/hQ4CIPeVMaUMndBwF+kwMksXvheRnIHLql8/FShcQ41SVHzY3afXgQys4k3WpaJOYPvlSAx
ljR4DhLm0JhWIg3IglfYTp2gd7sS9grQRN9+GjLa5hxXavGLJ6DWVSg7vYWTRSGByogm0Sa9h4GMq195YwJtiDpnAWVVHivKDTBw8yw4csHD0hCxn7VkoboK6QBBI9jj
+eNaaC9mYP9rkl84BF9tw2i4oLzESENfX3xtj2wUKEDKiCbRJr2HgYyrX3ljAm2IKbAWmvuvd8ilV1icDV9dy8BLGX1UQGGlSBs0L/OYhgklTGu3ghvlCYOZ80U7ddSl
WiozZBD53nvxqcPiINtO7cqIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17lKkOv1tpoGkegjZpOahEEIpHHPeDsh6+XOz1zDB850ZcKILqpViMAh92kTQwZ529
MKS9qjr8DhbiP98e3EH+SsqIJtEmvYeBjKtfeWMCbYg6Cy0VxXZenqBxkRlLe29KQeEKnkX4YftAfS7HQPHtlvUOzgVhr2GoovWyiZv7yByJscESQBuj93nozknI0ZC5
yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+/qK476G9VDG4IodOsSwJNXU49K9e5EKYcQmJffUrf9ZCHJYLdXEYCcJEEEwPiQI+NuPcqjj4KMfzKD264bGZmd
9eAhsbYpcvuVPp86ImPIqrHGbFZXraT+x8oatlEIJqv7rICpy6vrQuFpgCGDT3b17X1q+kzj1ljCgv3p1/3pwS5+NSNPc3P9ujIbdyeQBTreBEehDRu5tBQw9W4ARUw6
aE7tq/7wib4HT2wPH0lGOAJ5mUCE9S/oWA/UXCK8U5enNCH4rJdV/OkJe9vU0zdqnZmsuqL6lQq2Rh+X/W+b9cqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFz
/ftRmpGOfBINtgEt3ArOj0Zrvq4RiGD9XR8fLHApF1w3GoTeg5iR2AcMb4RSoGRs+UaZi5w/xQrMcnOMAGc9JyyxIv6RCIDGGu0TkZo0SvTOME33e6e1TCr6rznNWp7L
CJqQEctXf164rQaKB2wcOJVVYp8/yIukBGvPLOwo04R8trsGxbUD5dA+UtIyWE2P8irBFiq5/W4AZPCCvyETtRdaBhN59OBztKdEqNin52lGUqpUNe8Q4/WTm+cRfQkX
KKWCDtTSwL/NbI9YVYIv/0lXQ+GRYKordTkDtdaestB5BMIFRPGZ/oZOwygPBEfUwsc6TpcgBJYy/UwvWXMX91RLUwa2rymkJ1KB8TuoRHBtR72tobzyqEjMedAI8Lif
r9QsWLdQuzsj6jpaNSqQtR5gsHA9stndjJkvtKkbOIO8Kjycu14CCTTzXihWaTYKqmvt+9RJG29CVijnCj5p6jKZKKUW5XhDZ9NrPyOpABv9xSiIJEwYsF6cWxi0q4Mi
FRe8MsfaJ/3lhUEcM6pUCSuA5qC369hp3Yh7jiTowAHXXBAC6Vx2VUf6VLxt9KnJaq6RXpMkdhOCs5PZa7OpGuix1DERKhAVzmS7eoLsixOZF3EG1TvYOsmSsQGULznq
fqYO561r2b4meLoPn2AMcsa1omAuN7tugAFrz+M154u3+pVLi6r/cN5O+bS9us8DoLSMRgXAWDpD5MAJCsuWvr/P/F0SVf0SLj/NuNQ+fGQ+SxaBk0qG9B9pzubLYP92
fUgoSjZJ0mfLOvTfraoVzqyN31AZvu06PLFG+4zR/9Q3jRdYTEzTYQZe7o7yKjRVflmHgv0/Xs/9R7hHTn3Px6CgQLF+N9m4erX5R6ipBeKs0wAoZu8D0EYtW7hceMH+
85yBiGiInO8MlBueHOsEX8Aj8V60EYLqnE9Vg9aZO4E9pmM+AQubxtLx3XP1IwbG8wTg4MnPYNRzy/sa6yfoJyxBvbZGc+4odFDp1YqYou+FHOcwFzwhTqXeXM7xhSIU
bl4xPg643ANnn3EmekRHoXILjpckxD9y2j3EhJVZVgSIkwUEg4v96tuhO86cONYeySaLzDdAyDWGF8Jn8lEAlzivKdI2Qo73XQE/Qgs8ZAdNES3/oz3ZG3y0UEJh5fSf
+5WOexiqpmOiYKIzYiX0cn4Q7AfqG3z31KKNvrcNGKpIYYQlwiISLejsUvqCX21+N4BTssn2Z18FY1FkC7mP5GrJpHsioN39JlWxJ3VhxOSvc4akmV4vkdNCDjbaFWbR
yNciekSarizz+gAGwa+duxpB9NevwCx3b1Gxg4L01dohFh6YvV5h2k9FO/wGVc0lRW7iBTqm3qGpvReXH6urUvDxPR33mpkusJbQM4SIMVAt168FcGb56V6ZTIMlQJUo
pIT4FgSijqNFt69cMXFaC8qIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPvYmofxul3qzYpnJ42lgzFZ47iQ7nBaKh+iDx0aaXgHgD+gKf8d3h/nMSVAAkd7zTI
yogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKoGQh522mDkvWAEykxtJUjLyogm0Sa9h4GMq195YwJtiKlR4DSD3lXNlaYVFddT/8DKiCbRJr2HgYyrX3ljAm2I
3gRHoQ0bubQUMPVuAEVMOp232QK3gvaFq5nXKjibhYnJ8PgCLzYC/VqdgpdS9WsvaJEFPP1T4G9Ta3LUsfD7iNIjhPUODMVs/IQDPrkR3NXKiCbRJr2HgYyrX3ljAm2I
r1c+oB+tsltP04/RF5EClBpnA+yJ8xEpLGj6ZEGCzLbZB1RNJLDOyhv8yd1suqBKQ5Fy2Di1f0mpTAseOJpt09p8KaxIxCfwRJJPZaJ4EikQHTFkmTmQAYd7Un5pgxZU
i2Brb2P1bNYdqcrS0QfexN4ER6ENG7m0FDD1bgBFTDoNPuD/8geIbaBbqMR4cMkKZP44UTGS0lSBq4+N6Qvx8Kaa3dULqwAjJq5GD1eonckr7qZX6//ardjeGERThQkG
cjveAzO+/7U58YwS7JUaF4Uc5zAXPCFOpd5czvGFIhQv3LDdW2d4LJrahPI2i/Px+SSkItzYv1murxIBJ0Ad+2zVFar75CagUuaDiSXJzg5UxpQyd0HAX6TAySxe+F5G
UFcMrN2wuVtSYnoCCJUovCisPM4vWHVeoT+eBLF1ZeIIcYFqLD64vxb+DjXf6ZBrxVsXGMOQP1jgsB5wHwRFzB3xNFk3tNezh29P5W30qon2uzAflGXdSR4nP5/retPv
JnIY+53k2a+y2FQaRDoc5ts7XrCsThraVWqwWVxyrze2MDkmfcxoydmbjXXANtGjrILXHiZyOkc7Ta51JphsY31IKEo2SdJnyzr0362qFc6Cc7OVuHLWP3n1UfjkjOL0
Uw5XjMASTNuOuDdQLgltL3h+7q6YTvU95oNST/E0HoTKiCbRJr2HgYyrX3ljAm2InkPELMSQBI3KYVRngPExRs4wTfd7p7VMKvqvOc1anssImpARy1d/XritBooHbBw4
a7mBGiMYgEeqocGXiESYCxUXvDLH2if95YVBHDOqVAkDKsBl2hYE8RoxC3vzG1mM/1HfW/s9SyDCwR8+/8xDNaWCT0UYL9tZoNNRqctNws0xIqmIy1VtUXlQEiqP6rf1
GUnjBL5htQABe/EhEMqv8ZaQ5ok1rD2jnlRJy8CxKO70ba8q4Ioec+l3/OxQoldW+AAgZajUyXIcEJBTK6L9Qc0RufRW5boVfFR5t0EuYzo5ig9oGXx0mToVnq+Jp6yb
QMk08PU2rqVKkF3Y64R/sGhO7av+8Im+B09sDx9JRjiD/fltsM6GEV86zF7n7tQZpprd1QurACMmrkYPV6idyZb2XhAjMYBN5u/fOrs51LRL/EJBOjO5eE2cMdFSq4+4
aAneEQlA4p52Cckh9TZuS+QcCea9HYTVuheqP4K3WWnsm6QgG+Evpo2JgZJM0q28TazntDzpZp7xB8xtw7gHPsqIJtEmvYeBjKtfeWMCbYh5H24Cihayu6ZOI1RLHJB7
+oI/4T1qcyUjIGdq76uadW2aGZtJAW7/hBnchCAxhDjJ8PgCLzYC/VqdgpdS9Wsvyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+/K1K8YPhnkGDwPDAGy4ya2
juJDucFoqH6IPHRppeAeAHF4FmWGBChREE1xvbkkq5/KiCbRJr2HgYyrX3ljAm2IgRrInBgZD19HN9j5BZzno1/+JMQF8tPpxEp1hRfme5Zvy3eLpymXJAZYTOtu6FJ1
7Xo6kW/W3f4+4rV4FvdP8cqIJtEmvYeBjKtfeWMCbYiyE+El44KvDTcCPQQq3uEOSJwdnrpqIbKBhhntmvAfsVSd0D6ejAdCwdi7spWsr4VOLwfxrw7wfDBB3youa0bY
x5jZ8kFvTV4eNUYf1pBM4A1mJgNEioRCNz2EoNVMGX3pe63ksUGPLdD2LX2p2NW2LaqPkIWv91xHrFXSEw2IX42QzrD46TocVk7yxJKECDYt/sdTO9YDGG3LWyxHq+kF
gPqWAXrddDboDVic5ksdAfME4ODJz2DUc8v7Gusn6Cc2v7WBTB91D0AELKmasUyMwoMLSGqjvsD3e0psGi9R4mQOmX42tAo0GXVaafQdK6Iwoj3WUvEuMEQY5AFm2DEX
6tkKMqjDuFB6AVW0fn8FSpjH2TmsULwG6rQLKiUCUFZkDpl+NrQKNBl1Wmn0HSuiMKI91lLxLjBEGOQBZtgxF63ANzZfL0JQS4HdTazT/sxEg3WViYIzhFCpWgBMCsmn
ehqU/RsiveCoe4zfA2nZBXy2uwbFtQPl0D5S0jJYTY+sHWfJJsdEyCwhjfTtfajkczwSP7xYOf/jUOC6NiOlrXoalP0bIr3gqHuM3wNp2QV8trsGxbUD5dA+UtIyWE2P
zilpdbtv/nX0MSRs2ZKjtTr1j7+vzNEFtUj/71xmXIR6GpT9GyK94Kh7jN8DadkFfLa7BsW1A+XQPlLSMlhNj3ScTQSYkOQnXJhM8TsXPkWeXxMjZdqqFfLB4dLebk87
ehqU/RsiveCoe4zfA2nZBXy2uwbFtQPl0D5S0jJYTY+K2StNFLnGBpZyCQHbL8w3Ww+Erqn5vFK8eOGRKzDBRGk7Ti0yFT/PhF6DZ/Ty5xUVF7wyx9on/eWFQRwzqlQJ
CtQ/ipbaLhp3Emdy0R5aSDZ6Zm5BXDCIqIIK8DldFXDp9F3BL+09R2/LIFPpIP1mrrpmJsl9+1HJQVzeHhn9xt5Fb6NEEKN4ZB24Wue0Y3k0SrdA+cO+XiR8Nzc9Cf9O
bomYRt4imRitB36Eg0ga7VOnSXYlm9rWFpkroZ4t2ZmXmWTpl8guV5C0IVAd1NMO0B7U/QUqN2GeDPuQtfg7DbRPitmyAq516sxogUIJLFiAPNKa6BhT0CreN0YoDO4K
V8IdjG6WAFh3npcTSmn/VdSQfy9eaSUrRdRyOCDS744DqiWLLEE9/DGafiqNFrvXp7sg+lGqFJQp5uStXp9lXpXm6x1w/mBscG3yv176woYtqo+Qha/3XEesVdITDYhf
MFnvye7G5B9BPjubOa9rGRA0cRYQWHYQDQ3afcnMEhQmWWypthDbfU30U3ps0DW78wTg4MnPYNRzy/sa6yfoJ/+eYzXyacrayGcaw/mwa//SHe0BtRJRhOb75M/06LH9
72cnDLGCXm2170Qdw93kp1WenTDCmra84zjwxtBf2iHkkR2fh7tsFEruRd7sriOGWZvic3fQZ4/eLj8LYb7tbBYiOPAlky7IGdveF5LXW+XQ9oc7z1AzoG6bh9Xb1B9u
6iSDJDYdv12K6Gc0O76GlROskhZE2tnQbUIuQb9GP5VJV0PhkWCqK3U5A7XWnrLQtYJfSQ8PGe08Z43Slzlscr+u6sj7/01Y5CRYmq6/By7PzgzLSxrXPfn3ozobcl5M
HTmfdYSbaKVeeMXh96R53+rAJeJ1PxxlVYbBd0vPpCG3dqh1IL3fJ7NragoUoZcvT5vVAyEBraDCmrCH7htxRjcahN6DmJHYBwxvhFKgZGxTp0l2JZva1haZK6GeLdmZ
tGjIoNpp7BQP7Kke4J+qs5a9BosGr3pajxoYpi/7DelJ5Tq8Zx1zTjmaSNKuzsol2KYi8+Q2S4l8Hpn/TUcmMmy/+3QhWCaR0htFcQGGVqp+EOwH6ht899Sijb63DRiq
rJnIUp+6daRMWtVLk41c64NCAjNU17Jiy9s0i2TUkHh0ObT3j1ZlWsGblPwFhWqkr9QsWLdQuzsj6jpaNSqQtU6nKKtbSUs15igzG37zjfM7aRiHyyAhBTD0bKMRoFJ2
i1LfSHL7meCZLO9MHcLDPL/P/F0SVf0SLj/NuNQ+fGTYikPWyLptUvz6aA7afDc0H7qsns+3drobOr+zOqQIWzcnVG8fGLfziXifK1Obp1a/z/xdElX9Ei4/zbjUPnxk
wh8ceib41LiVTqXJ8QdpKDtpGIfLICEFMPRsoxGgUnY0L9QORpLO3dnyD3AoGjIBGFNNjWntikIRKxluogPwCfUzScAn/MLBl4JLApLGWIFLxx8cAyce+S5C0keg3otj
lElxNda0gbT6Ki+IGdg+9hhTTY1p7YpCESsZbqID8AlfCb1xGowBQQK5waeI+sUoO2kYh8sgIQUw9GyjEaBSdouVx5BpZgZzJJyl2Gs1AfsYU02Nae2KQhErGW6iA/AJ
Dx7EmTZqu/JlLjaPUFAuXkvHHxwDJx75LkLSR6Dei2O7v/p+y8wioa9+emlELHHJGFNNjWntikIRKxluogPwCcz9jnGrm0CzGA8gTq1iTtk7aRiHyyAhBTD0bKMRoFJ2
o/mqlwy0XqeuAAKt9mvmDgxgPFjJpEG/afkuVi56AgFJ8GXh26rvWrSK1X1CqgXupVnnu68LGZMn5jrT5JFMh23QNsmp+XK5Aor+YFzcP1OZF3EG1TvYOsmSsQGULznq
+nL6D8FishjbN4eqaykLxku3Vri+liEoGSD9vARQ7rJqrhay4gq7hsSMb6IB8RZR3Dvl2UwWs8UGRuHmdnMbE0NL3pDYCNd2/nB4usPKiFVngyeLfTVohu9EAzu70I58
IDMPaC3J1Si+R6jzSj/+u9rOGyZsI1Gj823nKtdPCvZa43zOUxFI0q+5a36QZKCwZpybsZrXNKq40Ho4H121fHy2uwbFtQPl0D5S0jJYTY/02n0BS1Jh7S0nSamh15e4
Om7nmn5VkvPfMjlGZ9uI3ufAfIvCERXvtTLZaT6qirbT6E5Nv8/9H8yn5zTB5EUwF8Mtad9FAmBDWvD2JdTR/xV5ECxGQ9AkfELIrWkEpWUMYDxYyaRBv2n5LlYuegIB
zuN02sK00v3yW8ipwPhfOpkOzFxaDfR36N6xd69vdoH8wd6Y7a9cEapX0K96FFHW8wTg4MnPYNRzy/sa6yfoJ/+eYzXyacrayGcaw/mwa/8g9keKryBZUTECjG2IL5cA
mHFuG+vnzJMBV/REA+ydfBy2ix4FwUzbMyaPn9APi9LCfzzfqevIE4pJo8iqr7jo0VpPB2fU0Peb4Dw7e11ZdQVAaYnzU01nb2xep1XnWhodDzvCjNT77i2NpjkAPOm8
H2SXqdCNUU1bE9TudIL7OTs+FcowHIPWZY/nMBcBQ14irDwyxGQu0fANTgmybZntb2c/FhwgFm76cayrLhJAP8+cxH87G4tuQiOYO54g89J0m4EEG9mVJ17dWE5OAOZ/
UYdBXCqRSISk3gHW4rpvl1DhScGQMisBMGbux7SOpXxheJ9IRFx6XeW0+6/0D7sOncxhybGbm41IXCy/t2uTwzs+FcowHIPWZY/nMBcBQ16xwmEtcPImN84if/0p/SR6
U5sfrIsuBQu+vYP36m19UBCo+ChGwmaMrIlD8ZxSSYJwYouYK1cSQoAyJnrbGpWxsL+l5ixmlP3W5K+q2vbiZzWSofj8WhNDWYVIvwEAltcIjpgx6oA9y3Rt+WffuzWN
Oz4VyjAcg9Zlj+cwFwFDXjND8vQzt7SPSUitjkEc58Ya4GA5CQIF7eHEJZNf2pVtEKj4KEbCZoysiUPxnFJJgsGrU6yRBMtDOjzHbk99nb10m4EEG9mVJ17dWE5OAOZ/
NWCwylNI/f82n5duGQOBrlBjqhObQrj76C14nS6j6Xq0ah3bjQWDS6/45tzlep7DWRcR/G8M4mq5Zr4+HDgmmVgF9GkqvI3T532KH4N1qB0VQut9iGGsiGExIMSkwCSp
LnCuiID3xJMB6jdkDBbgyEBV+WjpqJjCMAe/tOzGwrcS6+rNlYtfmm2dfIch8LwSE7ljj5TBR7PE/nppHl33kfeubT1NY+WcbifVjzBD2A9HbE8R0jHvFGkRAPbPyPGB
+jy+uVLO7P/S9Rj9eb3t+iwGeHMZIBq7x7CO9/hTJedp9x/TVikdNR+F1KSEHESYoyl3CZaFTaSPjcqO4UtRy0yR0wQ8Tx8aH+LJH8qtn1eQ6gL/C2xyi5a4TWEvdTpd
XrRdp7N7taUjSZwRPDNeedrJsV2I2e57Ry6qIjX+ZtWnYGwrtA1gqd79KwlPG4lF3tg36JZIjTN8D7VQ9R/VspNss9Cuj5M3gitJVXVNxZ5p9x/TVikdNR+F1KSEHESY
4zZDLt1vJlvjv/tdDo6vZmc8PEqC443YB5wHsuE5kzkYXwUFUK5l8xO+zmuxZFIMCAx7c7FK+3jtNkxkZTlIsDbV513lc3/eEEYp5LP+NBFJUzZxY2a6ArNLD3D1dmsa
Cr//AzVYWz0omU8ZPnMGJ6Ux8CDXSSmptXyrUVOAGfwOBP4XFWBudQ1ycW2VQE6/+XXQkgUyKNPK/REOg9/i//qwphVAF7URvS/m8mW4i560ouNgomzjPv4xDxjaN1sj
foLEl5WJkd/L1C3E83iDb7cIP05Ki5S+Xfb2JVkQvvWnr2LuqM+SIzvB3zE7xv7ePcLln0/+UEQh8oNs6DwdMHTqh/3se4enLlTpDFlH/qUhSPbQV3GDkoxJOSN61w2n
sTm07NUwEoEkkVHRGRuB6QZ04ezYrU7oTD1ZZ1LK//+Cpd3XQsOlINo0hYlmQ0HAVahJUgliMRUyZZH4sOfpcwG2pluJjlh1h4GMsQCglKMb02YJ93PZpsoWZxIbMny/
97RSH0WHudL7uXjKD9rid2phGdvm3YOZWhaka2EOg0WCtmkXihh0fDYLieB5jcIg60HU0YxQiAKv1pyA5L2x/YJLBgbw+OMRpkqsVZEdllK517tTNVAMplfz+cvhlnRd
amEZ2+bdg5laFqRrYQ6DRSQsebBULIi0f7Lm9iOEUDpNS6ZQn/3EBFjmKDfPhu3q52DH9FQnGuvAEf7XxzS108qIJtEmvYeBjKtfeWMCbYgoTSsTpr8+9n6cpuiGaY4p
WPhwY/5UmM4p5L2BfIfWmkdsTxHSMe8UaREA9s/I8YEpz41jYZgt7IKtAU/uReHc6kMkZ3Lq5ERp2HPxPzbxrARhg9IZizRFMSGUuA0e9IcmI8u53RhfV61/4IZh57M2
rZY+XdSkH4lY6omSSWNTV8qGAreB2bHy18C6e47KNRnBrwZZAbTiws17NmKj98u+xm1RYFBOCjrDYIAfpCyfjEaAwC8QC+1p0eETWnlFQ6o21edd5XN/3hBGKeSz/jQR
GF+YmtSZoTrOjZt84K8eEMqIJtEmvYeBjKtfeWMCbYgw/7o7cbYcsq4RNXcWtQPetpIvg8s5nR5sHudZNVeZ7T9pK7fYS7aY8716jXnD7dMPNG3hAen/DrT0s+tMr5LC
uZDQ5+hSUordlAPmzosF9FFVAH2U/F5RJ+5t3S5icYVpEe9B+IMMgNGFkdFTYOFZ8wBSbzG64J+YxKBPynkpoSidJqtT1R6+gdTiRpPojaR6E9EBAjPDutwdYiZmPqaY
NZgIQT6lYOnDvfO7a3rvI+GvAB9EeOdiIlQFpYU0J3ztOraLK7+vWcQ40D7padWL2T21jr2FgyaAyKQYcXUV9EmV3UcDeLGhA/7PNcP63UyIQVC7GTwrFXvPJ5n8bre5
yogm0Sa9h4GMq195YwJtiHRDKVZNP4lSwf13PICjvgMkCVI3QfLkZlhMZvFqxXcBzwnaGOhNScJ+4TY+Rh9d2Cs96lNrXpgxFHbv+ydKvBXKiCbRJr2HgYyrX3ljAm2I
RU7c4+AcsoCp8kKEqxqyMihjCialeFGfuGCGETt6jAQSS6uGc9h77/zxKbyuBiPOyogm0Sa9h4GMq195YwJtiNMhkZz2RNbOtgwPIO+diBy5z+T45eLB4BbkQucDhWbg
2nwprEjEJ/BEkk9longSKfvEMErrZ5unsZoWBPJ0oVJMkdMEPE8fGh/iyR/KrZ9XDgSHcWGmIYcbVzvC/yUmpX7mnTLeZ5tEzgvNqy0AW7VAjfzQ912b2gfKY11S1q4D
tf+YGAIm9WdQQ6VKwRhgB0zPIeLec4AISHAwMOl2qK/+8I2MrxZZsu2wkBm0NavdHcskiWWRcAwAB8VxdE6JLF+A7J0GvaqSHBMhcC8dtGUosV6IJrNh2Ga+hMpzoFOT
svLsoqeOuubblhHb0JtVtokkjRJf9T9BEGfQkHefDVH/sTtW1GcL8ju+MpBGYjwYXFA+JziGBpD8kgNLI3i0ZeLQ4Bw/cTSIV9+ePsJ5eJjKiCbRJr2HgYyrX3ljAm2I
+tMevWB4y1dyaRTdpuDe7pnlbEAOZQIDJXV2A/etOu56ijmp7TPsHk8rdG838NL6TazntDzpZp7xB8xtw7gHPk9AHUqNPiKMXd6TmqYHnDFwqoaxWdqCtHVnFFqvNXyn
Qga/g9FZJZ0jMTBc/9bggJekWncd6OGKl0oODEYrDUIVeWSGm3el+o9uSyJ8+pEdfshma5gZ3m5WUZsPRTH0123WhOYf8lFADwgxqMjK6VA4lnwY1nErI8uPz9gHpMgp
2tMwClSGZ+rpmgdLefTJqevxOxKR/2HUDToL1WB6dePtXnbedQQ+oyvRN90KRdOMiJv4UYoEDtlkxVkH3JNmYYjvt+9g7nQZfJp9HyYByM9ceFiExoXsjVm/fv/YbdkF
fqubin2dfEPTsZm+W7yVXVBEUDhk2Dzld0/iwGYN8+iI77fvYO50GXyafR8mAcjPvlwTEz9S1po9PUaS9imRVE1f1XO9UCIe/WV27Ypqa5q/5a76pRodlmEMKgS1X98+
iO+372DudBl8mn0fJgHIz1boi9OBSxlMMNUAYuM99gBmHDgKDuonLHrWh5gCw1I4CMe4ttXlKO1dfFgz3hYDMYjvt+9g7nQZfJp9HyYByM9W6IvTgUsZTDDVAGLjPfYA
8cmVV4k3I9619VsS2UXDoopVUwMUXs7qDKWTnyWf/wmI77fvYO50GXyafR8mAcjPVuiL04FLGUww1QBi4z32AIA0PpPhTKyMH697Xt8/3DCPG2B4Y/wR+yKHAvhL+Cpl
iO+372DudBl8mn0fJgHIz1boi9OBSxlMMNUAYuM99gDglpzKBlGPL+TR3YwA9Fq3wcIf0Xq5djjwbzgww6AFg4jvt+9g7nQZfJp9HyYByM9W6IvTgUsZTDDVAGLjPfYA
MhHrMbxMt5KerYcYAdYWuZkEGSEXKaoodkIUS2TLfwyI77fvYO50GXyafR8mAcjPVuiL04FLGUww1QBi4z32AHhc3Y9Ct9BSeoQoG+TIrLHYvPio/StgZOFFS3xD/sSc
iO+372DudBl8mn0fJgHIz1boi9OBSxlMMNUAYuM99gDOjRsIbFGgJOmMw56PLzD+/7RJ5A/bzTZycLeCQjU90ojvt+9g7nQZfJp9HyYByM/b/9NFco/jXbHiflWiSts+
Zhw4Cg7qJyx61oeYAsNSOH2wRieJd1QQBkDa8iMpwDeI77fvYO50GXyafR8mAcjP2//TRXKP412x4n5VokrbPvHJlVeJNyPetfVbEtlFw6J0+EfXDZag5FaBv15rg5oH
iO+372DudBl8mn0fJgHIz9v/00Vyj+NdseJ+VaJK2z6AND6T4UysjB+ve17fP9wwvpvVChahHCAhY/2hZGJl8Yjvt+9g7nQZfJp9HyYByM/b/9NFco/jXbHiflWiSts+
4JacygZRjy/k0d2MAPRat+7cE4h45rqBG5HiQkWZiYaI77fvYO50GXyafR8mAcjP2//TRXKP412x4n5VokrbPjIR6zG8TLeSnq2HGAHWFrlFRPnE0+fAaWvSpcNNAnIr
iO+372DudBl8mn0fJgHIz9v/00Vyj+NdseJ+VaJK2z54XN2PQrfQUnqEKBvkyKyxTK7xgS7m1A2vtEGCIreBGYjvt+9g7nQZfJp9HyYByM/b/9NFco/jXbHiflWiSts+
zo0bCGxRoCTpjMOejy8w/kuOar2z9V22MUCRAJMJVfSI77fvYO50GXyafR8mAcjPd9Z+tVkC7D+bXTzsJqPqNEE2GlQ082vNoSCLUj2rsEOzPxDfumxQdkY//rAxeBcq
a2KoULLq6hypwk0Raj1hjaxOx5vNz40/OLIovBExsiEJ3s/EKB9kDV/lGeqTBQcyXHe3IihnNt6iXfRJyWu4TByqi/W4OsfxCO8sCye2Rlwjy/r/0NqksMbBw6r16FtB
zLPVrqyoeXvtbFxnytfRoQKO4gc4GGYyfrah/dGVDd+KCzSldmBLaCquF3jtuogou/il5rpJsRGVof1G5ClwVdml7grUhnUSMSsZjcON72YzGF0/Y0f6/90A4ihb0ELD
Cs+bemYPefUdBgzoWZm3nCjBIxhqA4ljoodFlnmWH3WTBciGSAg5YGswbQBqSHk3nWMNnCLgt55q/BtsRxuV63tX8X7ae2aiup5kPpCFysKWY2ct18XFU1Bujr08Rtzg
bqUE2DjLiGZLZPSyqFYJIhyqi/W4OsfxCO8sCye2RlwrJcxi/7w926yQ1OYBH5RyzLPVrqyoeXvtbFxnytfRoehl3sA4TcqFMnR7RigbaK+KCzSldmBLaCquF3jtuogo
zhK5qGUxrOcu1zGeeyTBttbVbzW8kYeK8dQhs3BrSgczGF0/Y0f6/90A4ihb0ELDCs+bemYPefUdBgzoWZm3nCmig49lTVU0PIKfy5nInel64Mx+wYT8f1Wnxr75wPhp
nWMNnCLgt55q/BtsRxuV6z3Hq3zZGNWMB7zBEVjGonzIC1Il0xl8n1wUwHBXjZhwMI63Xv2pnthkdXuIlQA1PRyqi/W4OsfxCO8sCye2RlxzCPW+tnDgOblUzH4DqtZW
vWW0zlrdRR0oHBWz+iMkShjrwxAEBxPQCIuZeI0TRSeKCzSldmBLaCquF3jtuogokOifvVipHJTbxnuQiys6FkxuzVFYYd/3q+az+qcbP6YzGF0/Y0f6/90A4ihb0ELD
Cs+bemYPefUdBgzoWZm3nK3+tWaUTKfouCDpKfLJK/T6gs4cFRoQqIO1/6USFanRnWMNnCLgt55q/BtsRxuV61Cr/QBcLgotqmxsOgjLjf0x6o9UJm5ly7uIQKiy0A9x
ZWZawYFU6D99KBPmabCXrhyqi/W4OsfxCO8sCye2Rlwbrzxa67OQS1OiY2BG5O4pzLPVrqyoeXvtbFxnytfRoT1e2lvsUdURlYsglDwoKkCKCzSldmBLaCquF3jtuogo
0vMcCOUi/Q7Y3YvJI/1lUwNlVTL3jVsP5IXPfL1LQtozGF0/Y0f6/90A4ihb0ELDCs+bemYPefUdBgzoWZm3nCJifxtUm3WlhDE9aHgWLGnCO8zH2xjX5GA+Q5ZwvKJ4
nWMNnCLgt55q/BtsRxuV699uTvLZt29/INewFUApzc0pcQMGtxzrujk74VqroIXTyd7WElAuE3YZT0lQpl+0lRyqi/W4OsfxCO8sCye2RlxjZHFlPfycbG7Vz4c7lpwn
kmLdEUNEqKrPKHdXlwh8jGc02FCp1GXlEz4ytnzf6I2Csr9x9c98JZgJM75PSugDk7VbX3pjY2eP1T/APfjzapvFIuYR9aGNjhrvmyjgI5friEt0bzxxIL+02eX2H5Ew
tpBtrnD7HWwKeBej28173mf5Ryk8VJ/sXWDmvVzz2dfSdxS3mbkrCJEBYDQDbSu8zLPVrqyoeXvtbFxnytfRoXQLRn+8Dw+wuO+gwNrbLidSo2ZUfH2fQzOmFdVJFvzi
q16bTzQCybdUlPAOQmwbjPNX79aW59fBbfS+RmNyHERgczd1GQtMEvuyKGYcPXyx9Lug2+TdvjapVZC9h20rxWsoSz9v/i5yxQrA25LkCbdKs9ltzaplK7qR3naKFN4Q
maSqCZqJOiZ75/tZOhAPYbowitZCcQrPa+UP0SFS3DTOErmoZTGs5y7XMZ57JMG21tVvNbyRh4rx1CGzcGtKB6j9w1QSsWX/ToXozGIJLkfh7vdbp/VGIWrJvCmBgibJ
7qXbCwNzTG4DoEyKlNI+udaaAGmZkIliUhQFZB9smM2zIXrklMWLnXF8FRVRzHWbK5TivjNuJpbwi6O0qOC8fEIvsiuKy043oiCmebQAZYUyFuhwAG9QpZSwa1NnqIyD
XrsSePDsBh7vVQX5VT/nfGDSF0MR92jpH1JxOiYDZXaHIc9QrJiPwLvH4N+WdcKmxW6/HsCZLKWaNYAcvvlPIWFT1QaT6fxVi6rt+x9ns7jMVCalZmpGeTENrRTT3CFK
QyXTvScOYpYcni0kH7bKDVUFLI2iS/T1Cz02gHXyEEwn/Fx6KhIehIGWxwiF8yLJiXA0WBC8xEQCdhWVCg0vs2TfmkZz4U6vT5cMt4/ELw7glpzKBlGPL+TR3YwA9Fq3
jqYm4jIsQ+x9VReFZ9HyB915ruu0xtwCvxVUqQipo1uE8rbbicBKO1GdMlhTMy8A7HE/UfPo7WavMPLX1GxSduaBVdho2Vv3q1bwFtLHO7FANfcDeS6uu/8CyGTMny0V
YLLYgZrnoUHd1UOCfe3C3oaxeYrg74+r+V6cpotKhneNbHhuUFJOutkQCPzExFZ7b7+r9BGingpeOuUwolWMU10OOpKSIlxGlVz7XG8G4CMqQ+VU7VSCNklBlrXlZSmQ
cerzXs+a/G8fpOALa3xbUxPQ9Ge7miU8RJFtaqv+5aepminuUlCwt8d7cMchMDv9auCeHp0eqjyXYKZczgsF2cgyBsA+iLRk2bSbtkGzNGGvhKTabIx0JtKGKqiJz8o2
YYqGHDYFPoR4aw9COzuNwM8kRNRm5ZUa/YCRBOGj6CG/OfSRvNKbdweXQDj9UXRc+SzdnJcRj/iEVne6rGWBop09pVqkpLNQwkixjAPqRrmy0+o0Z9ab5t1zF674feeO
Cct/Vo5U8KlSiGTwHwuldVr+1optXfExfhpTywukv/Jtj5csJzPzfhRQf5/Ms58PRUulL+gIXnmDTZBPYwl56a9M39GzP9Y44muEF0spmxeCPD5vYVYUv5596zjyuchn
UMMTwYb6SNaYIRmECZKdQ6Qtlgvq5Hp/YwOX8NE5+nmycrSv2alQIkKjsDQKdHG02/bKtlshAIdjfLyduhFtRjp6uMp4xH9quZnxb2LyPcL7JeR6H6QFLzO40+N/CwvX
UwogEpXICSuAYgYsBI25PLv1KYSLvf0bnvV0iUvk/RFQq3d1ierFl25AmWFh02w1r0zf0bM/1jjia4QXSymbF4I8Pm9hVhS/nn3rOPK5yGemJ2NoBVzl5RHsS96BpNSW
pC2WC+rken9jA5fw0Tn6eYU8/qXn/MZv5R+KDWr25gnb9sq2WyEAh2N8vJ26EW1GOnq4ynjEf2q5mfFvYvI9wnt0laOSvJqFTUZs26AvyRcJAHvKjlRMfPEmRc4d4n3d
u/UphIu9/Rue9XSJS+T9EYpF7eMFD5QHaItDtxa4vvuvTN/Rsz/WOOJrhBdLKZsXgjw+b2FWFL+efes48rnIZ7sMqMyfp6bvv1E4M0XNDIukLZYL6uR6f2MDl/DROfp5
VuFl1VaHpigKv3B38GI5Y9v2yrZbIQCHY3y8nboRbUY6erjKeMR/armZ8W9i8j3CrrNEnFUEaXK6BdcvqFHGWRUx85CmNhx5EpTCWdEb7Oi79SmEi739G571dIlL5P0R
CTSGl+S5mbTKImR3+OhYK69M39GzP9Y44muEF0spmxeCPD5vYVYUv5596zjyuchnxYzw89pUeNBEzdfHRIWgjqQtlgvq5Hp/YwOX8NE5+nktrf2Tvr/D6QoBZj5iEb6v
2/bKtlshAIdjfLyduhFtRjp6uMp4xH9quZnxb2LyPcISlCdZv4smnryl0w6d6g7Qd6UveWk+p54IcIeu2BycoLv1KYSLvf0bnvV0iUvk/REtm6IYkF+yU4SHqYWdu7Be
r0zf0bM/1jjia4QXSymbF4I8Pm9hVhS/nn3rOPK5yGf5STR4oXC2wW/pnLj762LgpC2WC+rken9jA5fw0Tn6eUt8sOhG1yEpjjK4HE28CqTb9sq2WyEAh2N8vJ26EW1G
Onq4ynjEf2q5mfFvYvI9wo6REpJv6XDMTI8Nky76bYJzvWY4U+viHftCHtqpqj+4u/UphIu9/Rue9XSJS+T9EeFF8WuOZlOCO8xpNwlSCaGvTN/Rsz/WOOJrhBdLKZsX
gjw+b2FWFL+efes48rnIZ++S0ukPEHFNtScluxNMNRKkLZYL6uR6f2MDl/DROfp5nDXn6O94BEclEn4vl6+93tv2yrZbIQCHY3y8nboRbUY6erjKeMR/armZ8W9i8j3C
+90iiKAzsPFxjOXLyqS70Q8kCktoPk2Yyakr8jwvfLW79SmEi739G571dIlL5P0RNevTe52dnx5Z06ronZY6cK9M39GzP9Y44muEF0spmxeCPD5vYVYUv5596zjyuchn
8E9NB2ozSBdqsOOVOZsoWaQtlgvq5Hp/YwOX8NE5+nm/fAL5IkzoKOvmH+HP36Iv2/bKtlshAIdjfLyduhFtRjp6uMp4xH9quZnxb2LyPcL73SKIoDOw8XGM5cvKpLvR
c71mOFPr4h37Qh7aqao/uLv1KYSLvf0bnvV0iUvk/RGQm8nRZDoHUrL4roHctQKBr0zf0bM/1jjia4QXSymbF4I8Pm9hVhS/nn3rOPK5yGdQwxPBhvpI1pghGYQJkp1D
pC2WC+rken9jA5fw0Tn6edHLTDNb7oBH6UuUodoeaGfb9sq2WyEAh2N8vJ26EW1GOnq4ynjEf2q5mfFvYvI9wvsl5HofpAUvM7jT438LC9d3pS95aT6nnghwh67YHJyg
lAdBphtu9B/U+31q/ER47LriYh+rYxkqZq3q8C+GjiaI77fvYO50GXyafR8mAcjPj3XIukLNJKiErLWmtof/2td/CZq8VSkShlB9gLLMBLrhfIViotqwhXYxW4oO7JfT
0p3GJ+vojM3HcGnOAYd0m5W2f3SkAPTfZlUpulc4w6qsTsebzc+NPziyKLwRMbIhCd7PxCgfZA1f5RnqkwUHMm4thwY+KMBbg1AHLr9CYdakLZYL6uR6f2MDl/DROfp5
hTz+pef8xm/lH4oNavbmCdv2yrZbIQCHY3y8nboRbUaIguZtZjG0gbEe55qFZgFvINDCmURftuqRP4/wK49sRd+TeTv7HUuyZKCPaWinZ/e79SmEi739G571dIlL5P0R
UVBsDuZXM2oOVJmgC/sCuPetSo46JNIh2FMgyDkdWK6waeWtLlj8bJve8ql1u7EjzvZ00Z/wbiQnZtOAwDFOxIJLBgbw+OMRpkqsVZEdllJ+lGIGHWl10VqSrmofjPrK
BXPwLws+qCjn53tpPjinDrniZSs2iCi7ZeesRoIQJFSbs5SnKqv2qN9897bs7HoClAdBphtu9B/U+31q/ER47JWlUrHciYtell3CmWzYIndD5+VEGNCg7Q+UTe4hT5m6
WeHkYSVv/YWlhkhNsDolmNO5Bw94Adky7FjxdBZXIduQ8xxgnqIAJkMM4Lq9agZrYmamzvsbbEXV+A4ycb9XF/N32f4VYmoOvIeX0kfMkD5+MOOPJIBBKC/oTL6kqPk/
Ucsdv9QKuTyMiDh7CnhRqlnh5GElb/2FpYZITbA6JZiIL2Qrllzq7oZ1+3/zGlcxbnQ1JCQVFySJH7HBtixhgAQXK2YtWpg8DNDYn7sjSymfwvD/VwasbXrlfhyvBFQK
Acs2jVC8wcWHV56OheD1S0biasi91fJzfL7jHYFyfQ0Oc6LQWKYaNMe4k1ewXbcqK+ynFg16FuLaPMd/K8kpjS+21czxocYVpIimVAPrhKcpJiKsbEV2MpnLioBYJgDM
RzyuOaZp7cBNy9MgIwOWVwZZL4JpkPNDCeBhZ4t19lxsd9rrFHh24Z17Fqfj18VEaUK6QNVwqqyFACQOyf6Foca2pJ3g04WHIMlIJj/QeV4wKW2u5lh/DiNlE6eGaKLx
8hzkm/cA9HRL66O/qFHDTuJJ0wD4+5wSgJ0WqALdtDTHOucAxdE18YYfdb+lLZsAEp+e4vRsQquPBMHPirEKESsZz4w7OdXltnDZs+w4Zi3HRNPteYh6ngCYCOnDZNsP
0e7R5B3wOr48yiY2Mw6Ih+nu93NslJN0quT9FiMD8u4zon/pH5UlF29wr/WSArX3zVOQgroPPZSc5M+8vafUaYWrIFcfhrjNksZC089Is+V/EtaR/hyfuxj2CHDqGvmV
TJHTBDxPHxof4skfyq2fV3B9cAEWRn6hSLCTdi1z61+YQH+IJq7c3T7tA2iFcEDoVL/BrS1+IfmWhA8Qnucvz2sJZ9opP98H39UXoT6bKMnscViM8CTU9rHXhg1j95Ae
BmSMXvO7PoPY5FKgSy7gzqdB1KV9HhSx2fZmQRbmqESWDHg+NTw8BZpkxWRRNJHh+O+6Uja0DW3I/RLNKCvmPkOcuQB6xJQ1Ej3Dl7Ua/buogSQ4fbq1Jvd16HzQuw1Q
hHC6BVXmqgfT10idaKjnO6QLueb1eXccRYIZgRLI4HMQPefhLttpp4JvBefZQdUvLd0GtWF3SyqiItIaQhneXMmoJ64B0z0q0Qo6PsILL9RCLf0kpPRiMEci3OfmIUMK
yzar2rOeLj+T1gLJ5bS8N8a7LBSVuedWe+dSUqYFf7klG61hEgSldOiNdkpNFmEpk3c7NSvAd0yT6m2MZQLIObPE71fXEwGsnuJhVAocBhtA2OCHcce5DOGxweC7sovi
jrSKCqvS0YPzc2ihEW3qfoPx3JXMtWpuvKerxTUXbKOTdzs1K8B3TJPqbYxlAsg5ePqdhBAfrZJTapDvO89AB9/WLWtsBHgR5EYA6GMwTQjOaEdiNitYss7kQelk9ERe
8/gXwFlJfsPFgSBPiM8KpJgY+8jqnoMHNs/EVGaISxYGZIxe87s+g9jkUqBLLuDOJO59PffikhKc5wkPmP9DinhYAerMFi+knuGL5F+LlYl9Gm0/lcAvCt3Bl3G0Jp9m
q4n1ykMx/UgCHnJ1yalNgT87zyqR7BVFY7OfLEJl7+yoUIJ3uW4nGuVV7J156k+WR+f+Ql1rZhqjdm+V/vvTi89Z/RHB5c/ovOPZcNyhWor477pSNrQNbcj9Es0oK+Y+
QLHJ3Go+LlpjwXdxQa2KHQYEWKew4oorhoRSVGtr/xSkLZYL6uR6f2MDl/DROfp5hTz+pef8xm/lH4oNavbmCdv2yrZbIQCHY3y8nboRbUYJ7uqINAlxTNQwVdQNME0R
C1+ku/evEBzSK7+up8pTMJ0VQ7IaC7JEcGjMr88zH5Yb02YJ93PZpsoWZxIbMny/ejb+BXI2IFM7L/hx8D5hhAHE7xfIMKKDCpigK7+ZtPAEbOSu6bAZtBeUewmv0XD4
TUumUJ/9xARY5ig3z4bt6qdOVTyjAt0ziXHuykvcWR7Rxw8HqBS/6nhK9j8Dggr9CZLvqFnaYmytTOIi3F5P97Pqzge+g22Bp+dJaQJvBsDHvX+94cwjquOItOE/SLgs
KGK31Tkt1AHhqWq4/Fo/QoKl3ddCw6Ug2jSFiWZDQcBwyXpHr9liR1lLGX8/mvOeAhMr0ydlJjoIpojAZHq9tahPbh36LnS/oHJbkYg+Fx9Zyxs765Yl5pBuS3jSoMzS
U7STCO4qa2vS9NtKbzQrIMBxQBNES/U0OWbKWhwjZAfgFdd98i1+l6eWkLsbMptoZz9KwALhkEgKYIHHZR3Z69PeNRHwz3Ge0CBXOIRshSVR167TDTxyn1P5j13g13U/
Hjmas67PMNSXTU9VCJWmKmgHuK0mpGyLyLu/nTn72cecvzZNyxjg0sHeUiskGIkiB9wI0PUYksOZAS/FyvJ5OPsEZ+0iC4/92VOZfJbpTRYww6gJn4ytZNrA3AU/W50H
Udeu0w08cp9T+Y9d4Nd1P6/7B1BKuDupPT3LfPl86iiqJW+kG0ZGCRsM4llWbzV3UF1OXVfrF1t9Vmlu8Xs5eIK0xeQpcFWw+mBkMZI+N3JGVnYp5INQQ1rsaqEML87X
cX61fywPe2MvhlMyjb7PWzDh7H4GdlJD0kHbx5D5aVZfOENAw/5L/K/Wo8W/jZH2fP0ufS1/d+Ua92j5I/Vgq7aDsAtaQrUE4Nsa2AiIEIKxAYA9aoWHeA8YYsYfBk9e
IZ9iNbMLZG7R0MHj60xUU/5+hvjJtIlo86oVHNIhG4qMVk5iqZ4IVxVyZQhH+mE2XsSi4ZoQ96e0rIDTZiOPMoFIoJmuPfcnt+LYAPnEUDe65b/At7yQ7khThQd628z3
YD55elXoNVieDwYr2cnWiAJnSuw/vV1bKxVDZuULvNICUN52xnIgsllSngDLXnoAyX30krz0fEHwro2kqotauwEsCCY+4J/qk2llKXx3bMehFn8VIGbOtHDSfkfGsrei
nSSqVw8/wHqSonyLA9/sWLmQ0OfoUlKK3ZQD5s6LBfSG7m+SxiZUcxLt6UrQMTp62/bKtlshAIdjfLyduhFtRreHNYype4HbtYBYUPE9cE8KGxN7ng1GKWM0I4vUXfFN
ogADLblqyaL3KKB8o9hsodmMHL0DlafbNCJUaaFG9f4bJ9+EdVZVAnkruDzZuQE8jDZ6GKd9wnL0BoJfuM4JtKLmkYp5J1p8qO2tSdKwoNT3zBsUpqubA/RnFfO6SJAt
F0sOrOuse3pwx7lzFW2FNg1bROZ7ngw8MKU4njCC0W1nsyRX/H6fHyEVqlh06TA5jAxm5njcazN/RpTRaRP6EXbsnVcPsY2YVfGQ1BDCHlyLmwQkOyNIbKzPAJcxrWQu
BR8OSF1u5xKm+kYWq8kQfJUl2fJT8Ot7wRMN2b+G/5tQ7oi0osY8sDnJDwphQ+0l+J9h+KovGBMCYQa/Mj5O95Jj3LU7Coe40ABtYb4/n8NH6xOxSuYx0DATadgRE2i2
gBUXChQW4jk9V/40iULYjeYzSs/ieTzG8GBr+/DEITlRovCvkF0Pm9LnK6U/f57TQnO+TaWdJQ/PopI88CFP2+IePStPGhnptG5vwBOv6+a0NwOJ0T6HyX1RKvRK2/9t
4dldRT+0hYNpzp4HLg4JbadltD57AOFfUneXTvt9vJpo27rcbLaRRBTI5nNxPPkkuRQVGJXPHHVq9MHPz047SKRpOoX4B5JKjMq2GpUUOYSWXE4b2jIPP8igXhMLv0kR
smRIpnrgoI5Mvz6liOwWSS8pO6Uo138toTqLqthL1E7ppv26v8izE8cElbzefdRGbL+2nC9d4o8GcZGMNDAOo8ji3rGPP2kBW9NPG1+mwIXNzqr26LBZADP7KUNUK0Wy
5kKZyKMyc/F5jPUA7A4P7N73PWqsTBnhaWhDWcrifYCTtYeqxTIsyfvgtsDFIRripdFb3QU1zYd+ZoVcEpqceOO1HvdGPoP4dMYCtIC2S+MR/Ie8DbVlf9mTQ1u2rVJ9
uIaUOdHlU5RPvdH65BIVB0YJvE+Y+H7SN2Ct2sZ0flMh7zTZnG6Nz8izfLltCBGEqA95FKKKIFIus0zov+gm9mqIrHj3in6saN6Tbyepj5wko9HGnNC8CWItqYFFjby6
lCdSGvVngX1auxAGHA1XwJ7tTAkvdCBkWZPOxGc1VKmb2BNh55TQk+b8gwIF7NFpsU0r9/m66+kKrukNwKD7GgTqs7Y9bgT5F/79Km+rkEG8eMDU3kwq8F6AsCz++QZz
IJRJ8HtbnyyNvrQUxQ/rVr2GaIuIRFPSndE8P1sFm3zR37qdzHA/b9I3x6f/Xfm+uvSTHv7pZhumcyKpnWVpssrvtEHogS2pU5DYQ0Eey3FXSq2xzShHtfTptNGC6v+Z
EcGUFRbya9Xqy/Xs2H+2L+XViEHhbuAwiyU1Wo31MLupH0IP5hFhXsU3fKF4ag7g1NmhPqDRLNcGg+OzsAiVPhRiwHZJEJ1ypqqKgExMB/bNOjx2NWUzsHbv9u4rB9g4
+J9h+KovGBMCYQa/Mj5O9yrh0nbEaWl2E99qppGlyDJEIdZ2UMDZ7e5J6dTqp8X8HQ87wozU++4tjaY5ADzpvCgpqXE9q8D346eoFR97BawQiSzkvh5Gw/r3o4FAFGHB
I6hXTUvv6KBrCduTj7NNhuWqxgyPLqgXgLVpMHIq56FaQkdwA0sJiEf65KBf0YiYqlAti59YtJbRfNdVwFsq3s9YWInS4C5SzEaHVNuYCSIHAIezRuR6FcRxHVKJVLYk
jnhxsY7ZXzciPv5X4LFVFzs+FcowHIPWZY/nMBcBQ1597ZlcT+27vQTj3T377xOrviRus812Yn7eaN5QLUlfMZCXtHUbvcnUrHQDnnoZso7yHOlOaXcInjx0d/rBtWQl
2RSRGFSm7XHFhiZdlmAk7e9ioAvr6tftESnMX4cgPZdTmx+siy4FC769g/fqbX1Qo0NLXFlLfOh0zOdD7qaDGNO+wN3X6/KSPzo09k0vAhjpDwEEZvyPjqh4KSNVbSCo
vpP4kO1fx6PUz0G/FZb9XPCD5FNglprGT3JDJgCOeRsoyf5JULeMMukzOzQE2armkJe0dRu9ydSsdAOeehmyjqjSA3q+aADcI4rcxnTBTU7ZFJEYVKbtccWGJl2WYCTt
RjIhCO1KiriYlWVHMyQDiFObH6yLLgULvr2D9+ptfVBNbAgsB9nwqY1AEwyN50/no7TjCPcBdlGJSWK8Ya6qkzgFy7p2AZ9iO7hMJgaPzEATjGXnw8lQKbh9zZRldoMn
6Q8BBGb8j46oeCkjVW0gqL6T+JDtX8ej1M9BvxWW/VzQrxMUr/kGF2F3DZq9GrT3OQn+z27saTsf5/vBGJysxhsJcBqADRhl9Q5U1AO8e76+JG6zzXZift5o3lAtSV8x
kJe0dRu9ydSsdAOeehmyjnklAfibHXHrdsd3/hNPr7f4n2H4qi8YEwJhBr8yPk73X+FCdPtWVSUCwQ5APVzJ06ajoYxS0YRlvFOXimZ7ehgpCDcrAjYtmlaeyff0kPr8
AmEuCkHvxDkkAzGEXUHK7x82vi8OBFHtPcRiBOOrWsC+k/iQ7V/Ho9TPQb8Vlv1cX0/kq8uhXVo6ScWgF0TZyMtNAprDKFZOrSrNBnXaZRtew0ssq4VE8J0AKSTLcrvJ
2tpr/kifjMXfc/z9WExT15YYDit/xCmNY1fCbrQ8Tzf50yjg3JvUFdGSIDz9AKbnxJgT0pNCgmeSk1QS4wGXgfgwzH92yJ1yY96Zs7RW7QQyyfddVqfvmGojP4PrP+xC
32dn6QvycyTFS8gFC08DoCgwldlyIJg5Qz8/WU42V0Dww8Di5tSAZZkUZtkcCk060gu+0siZgpup1A2MoJfBZeByTThi14TxdAVxUn68Hppz85KGOCdgMGccuMhJHaqR
gX4ZSycEAfyUqd5UH8/+XV74WJSlUWNeQHlUHp4liqAM7gE7AGYFG4Yb8pAFf2DmefroLDhNowUsfK4GDEWja5TxTY9+VSAtep+PYBr1toIWovqjNzfwVrXx/La/Fkz3
UAaz+RuWwlgjbYR9bWYshG9nPxYcIBZu+nGsqy4SQD+QYhLJKCTHrYyrGGG/X6xNiTKXzDds5jGoH+lxuB+/IB0PO8KM1PvuLY2mOQA86byvGweLzYgn4KKUWTFHwOkH
m9gTYeeU0JPm/IMCBezRaRxOrdXUxq0mJ4K+s7B72YtPWAnBmKQuumFeIhGCajYeJyR16wcxiTMWFzm+rmBjYkaVIopWGvF9w8pYObcyg4MQiSzkvh5Gw/r3o4FAFGHB
4C68iIvmUgCxPUO6L+/Vs0qtCOfLHeq2Q+VSonDvxUyVJdnyU/Dre8ETDdm/hv+bHSAYeM2NrwqgQ1fiA9WjtlgF9GkqvI3T532KH4N1qB0jqFdNS+/ooGsJ25OPs02G
gwxvXRtSU2m15SluvHUAgzkJ/s9u7Gk7H+f7wRicrMbeFvXqaE2C3jSHxJjP5QpxVdzY3EiwwpZ9Sopd9kQ/pEYJvE+Y+H7SN2Ct2sZ0flO70LE+3zI7pdXwa3n1DvjP
WAX0aSq8jdPnfYofg3WoHeLI3jeI14W8cGWZxQYdSb6OaBNaNCECDVqj1jbqG8SfWAX0aSq8jdPnfYofg3WoHSOoV01L7+igawnbk4+zTYYOTJOdOE9YYzho504Cm7hM
OQn+z27saTsf5/vBGJysxu3XsZtTCVHJ0AWd7HJzLsVV3NjcSLDCln1Kil32RD+ksNrRM7pVU+Emssz3d1SflEld+teYumRIBPsElUMeqzR3K9FwusBR6RqbL2CQ0sTx
XFf3lnOlleeYi4vKZiy6K1gF9GkqvI3T532KH4N1qB3iyN43iNeFvHBlmcUGHUm+e5vuWQDgXqv3Xe9jHZ33bmuOQEBPgr0W7RC39cz56aKc6qdgiyRCL2kN8w0PhI0a
WAX0aSq8jdPnfYofg3WoHRVC632IYayIYTEgxKTAJKkucK6IgPfEkwHqN2QMFuDI5XfN42XVmXs04BAlOB50AZUO8R0y7/A4NeaU+32ASpE7PhXKMByD1mWP5zAXAUNe
v1udl9kjFDYudYwzbkr/G3SbgQQb2ZUnXt1YTk4A5n9N34nIA7DNyoi6052WXcOCPiNM1j5TB1kmTEVmEWdtOM3OqvbosFkAM/spQ1QrRbLb4wtfY6Jqq9ulLr9kLH69
pKzo8TF1jr4G1BoKtRb9p97YN+iWSI0zfA+1UPUf1bIAtjW3m2rtRD88YdozTcLJfsobjR2KvEY235srnL0HJYvKvqUAxMn1Yx/4GLU9PJUeRCgeXll+yWw0PYTf50uB
SVdD4ZFgqit1OQO11p6y0D8VU+CYr47dMnmF1Nyiq8dEx7SDuyF0S5IAc1wGiFcJIiycjjkTTbu0pW4V5MCC9Hy2uwbFtQPl0D5S0jJYTY8erSrqhA6LNbw6CjHoFhKS
6fe9MSJDPAhMU0akxHkUOTVSt+CSNRgdLFBYFmIZbFzYikPWyLptUvz6aA7afDc0q3J1SjMH1k4FLkVcmJSM3RwGM91Je7ndQoJOhBSVO+ctqo+Qha/3XEesVdITDYhf
eH/tIJ0OlQ2MpnXPoVJAwZB/keYmgETpbFXygYEtO2oiLJyOORNNu7SlbhXkwIL0fLa7BsW1A+XQPlLSMlhNjxSHpRaErirurfF1FNRgdLq+k/iQ7V/Ho9TPQb8Vlv1c
DsqYdBXv3mMn7scrRWeHDSVAhBR+E1z0Df2sfOJIOu4LoDmqlfjNoP1jM/eiYw7SHHFmLwr4eHi8nGNaFJfXE8pnqJlZ3Ft3skgaHMZe2p/2LcJmvrU7s9KH4nTLit/T
Cgy0NKkAjaL1LnsSPycgeSocHGKmvc8SwR0BUYWpiI0woj3WUvEuMEQY5AFm2DEXFB+OiPSYyE55etxBaeNGbBxZ0c9jEHXy4ySPUSaCHYUgNrZXNU955Pi6+BGae9Ww
b1OBWBQtoHE3axP0T1C61/jbgiUqlrA5YtkrHcOd8EghoYLzsBKAHDg8GFjNFAvxAxzkFJ3Vk9enLz4HzTuRfjnGkZnXMusnRIX7L8CcMqBHbE8R0jHvFGkRAPbPyPGB
qR9CD+YRYV7FN3yheGoO4PME4ODJz2DUc8v7Gusn6Cc1Tba0boXaSD2kgtA8983m+LAAYZ2SpYAdz/7rsgRCMJJ4GrscHaa788EgkEzXRnCy/apfKYtudsu6kQynVd7D
9HG8HfrOzrxBd0aOFH9hLhxxZi8K+Hh4vJxjWhSX1xPAdjE4r/yylCgkWJyMQFUI4DVR62C6aIB2Klc/IePDTXyHPixWIgAWOGUBec/OeZi1GE0b6JLm4hSzDp96ruQU
pKzo8TF1jr4G1BoKtRb9p97YN+iWSI0zfA+1UPUf1bKtRAZyrZoqIcbb1g2SqLcuNFg+Pie9rNSczHHrNnqTZd8ctBV9iAOJmsnxuiIIJObVw+WofNBXAcQxKjCDqyex
GUnjBL5htQABe/EhEMqv8SVqm4W4iUIAf6opdGDLctRGCbxPmPh+0jdgrdrGdH5TIDMPaC3J1Si+R6jzSj/+uz+rl30tmBgXrwVCsnyrrCEoVHIKMbS+apsVZ6zCe/um
SMi1WcNO9IU7Dx/SR9IPMhlJ4wS+YbUAAXvxIRDKr/G5mnEt8H6OPI0rX4aEiyL7zc6q9uiwWQAz+ylDVCtFsiAzD2gtydUovkeo80o//rsk16aj0rIWF2UWM1FHODpv
zRqFSenvVk0sY5jJJpVNhOWhLAdP/Zbp4vm7mPfI+fA5ig9oGXx0mToVnq+Jp6ybutKhc8+LyyWns+eG8vpKqUNQjGq8q1uR98i5cVJRU6FgI1gIhLNFor+KrP18O//W
dKONTzeKN/btwbLN5HrJSMqIJtEmvYeBjKtfeWMCbYgKtLws2m9Mjoku0HK3Fkm/lmZnVgmA8s9Dh5xMlj05uUdsTxHSMe8UaREA9s/I8YGBQUqdOoN0MhXxvU6NcXE2
fsobjR2KvEY235srnL0HJRBL9mFYvXCJjYl0M6lfezq/0pVfg2YoOAJHnnNGQ9B58wTg4MnPYNRzy/sa6yfoJ77kULT3zoUs1c9KA5UJw0GqMQbLTp43Mkw1DhNI++it
OYVsiatft+/31CXedmMNyBKEa2Ac2QN/Kr70Jr2uraEzxDlvZddknEwrcmFaq8EKrsQ/aeJOH6AvDNRKocmgC0lXQ+GRYKordTkDtdaestCykZP8suwbBEQWnuL2Zkrr
kQbEJeiz8a5Su6JLfydyXwq0vCzab0yOiS7QcrcWSb+PsK/wN45TbsVINR5bLNxiCXegWUHQf53gcMk0FUjRMWBGftxdlxIHtuizMMA8vyS0HfdueVTe5CC95ydSzFUh
utKhc8+LyyWns+eG8vpKqZCXtHUbvcnUrHQDnnoZso6BdEsGutJO70tMDz38PjYzxqpDgFqymu6ZCFhJ/bIRInyHPixWIgAWOGUBec/OeZiCFS8moB87mw7nU//gWrJl
umfcrKIXNsuMm3K+5kq4QUTHtIO7IXRLkgBzXAaIVwmadXTYIk6kcqeOXYRtqz63l/f0pxG0tL91ifOD9P338IJC2K8A+N8Bmwn2fb8A6aUPHO+bex6ghgxwpWbPVlJr
SVdD4ZFgqit1OQO11p6y0EAKBUK1brTy0PgLNIUJ/4Cxe9J9wbER5mmniAdaHYDVmnV02CJOpHKnjl2Ebas+t4+wr/A3jlNuxUg1Hlss3GIysJ25GTPKWsu5Kgw5yOCn
IrpITs4eavTHoYKwdprNELQd9255VN7kIL3nJ1LMVSEr74YghVdYOP30D+X2kcsn6XJ8OjKuZFnzOascrhY3iyyOgBnJeXwZQMCFs13/pW7ZLLGiyuxqyjDJRhKHgFPH
Uw5XjMASTNuOuDdQLgltL1yk7Sx6zxZYFWHn7Mz6T7rKiCbRJr2HgYyrX3ljAm2I0yGRnPZE1s62DA8g752IHL7Mbe8/j+Ht4dB91ap/2NpcgDog3tor3qUWo8jtdp5m
9Q7OBWGvYaii9bKJm/vIHPDALGczL/vY+sehpiDbKv7jjZyS1WBUX7rskkI7heHHia9fmNFgGjI/5LT99C91GsBLGX1UQGGlSBs0L/OYhgl89ysXk7A1qwDShe0ZKOOh
AIwHIyopurEKLePQsFbPvA2ML/eOYKfyOTM4wQe9nijeBEehDRu5tBQw9W4ARUw6DT7g//IHiG2gW6jEeHDJCmW/FIR1KBz42cBnc0HGyHsU4Cct5o0X9iaR+3u1mRYA
jwKb2xqzyN3JX/aaM1GF9MqIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0izjVrB7g80lD6Qd9W0lAUPX2HG7SxsAAn3nrf4KkXttcFGzJa9OWj+TQGQMtaNYeU
MetL3c2s01pfQJaS46LnesqIJtEmvYeBjKtfeWMCbYg6ZwFlVR4ryg0wcPMsOHLBj2GUcBMp2/liOgoQkvqJrbZy670R9qS0xyKBPV/qcM5z1Ofhdz2WoRv8kOx+BfGQ
yogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKp49kVNwvVhJPMyLFcZvXHgMSWKQH1CD+ja6FJ1FBewYlzZHkH5ksIEsx+SDct/K+PWbHX+sO+s26xbh9z4hsQc
yogm0Sa9h4GMq195YwJtiFBXDKzdsLlbUmJ6AgiVKLzEYfnR4RVDweW5WyzLPRt6wJ1/ts45Z/Ut+Y5yeQl3s+9TpxqP+ai4K3t7DIuL6gpjiyjfzVTPXrFbZ99I+uLJ
cgcuqXz8VKFxDjVJUfNjdp9eBDKziTdalok5g++VIDEA4AEl4pNNCx46HLNELETDuFF+e6TVrsoC82ybZql/8CJOI697b7CDHLEVyYSoyRnKiCbRJr2HgYyrX3ljAm2I
9rswH5Rl3UkeJz+f63rT7+orjvob1UMbgih06xLAk1cN8baeF+fzGrG2SNdre2qWcBbL1L5ZFa/I1DMoXY/A/wgsYLG4wUzH3UZZqskV1+xPQB1KjT4ijF3ek5qmB5wx
fTaaweHIYBzJm9VObDkLB1xjBTmwfM5MLdAhMd/LKPNyC46XJMQ/cto9xISVWVYE6FLNqIRc5wXKWdgn6DybdcqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOej
CfNcbnQ8eC8VC3A/6mcJ8Q7WxWpKOlTXm64evPTKs9gCDs/CBCupkkKuyYlwBRu3oB1H7eess8hzaBA0sl1vHMqIJtEmvYeBjKtfeWMCbYg6Cy0VxXZenqBxkRlLe29K
dCzYttXyKsMnnU2pzw8NgzSTHJuylT7x5N5x/ctiPigppKrFq7TF7v8IP4QzYF/2yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUYh1/FO5Da3rsrLoZ+FIpuO
TX90VAj5s2hN0DcK1cpi9OA9QX7IvxriU2pIPEiZKg3eBCDeb6edJLK2ikueWrxq+6yAqcur60LhaYAhg0929ca1omAuN7tugAFrz+M154vVSBTFAiG6HSViOzGLHd9C
2ztesKxOGtpVarBZXHKvN1n7bjcELL8gArzlDtFSZ9jKiCbRJr2HgYyrX3ljAm2Ig3EXTn58wwiGNPL7MS7tex0QxInfO9/I+uiLMBfqD9SsxKHmM3aE5Q+a0eaQPJKM
KKWCDtTSwL/NbI9YVYIv/y2qj5CFr/dcR6xV0hMNiF9n/d5WXoO4O3zkf+2jc9BheIJSTMxgJn4+DLS+j60TU5f39KcRtLS/dYnzg/T99/CQD9zpid5MwMawn4t+Ynf+
kngauxwdprvzwSCQTNdGcBUXvDLH2if95YVBHDOqVAmWYwXAj8HBupltqceN/Ilt11wQAulcdlVH+lS8bfSpyZDszA2YFzwuvKi24QS/2FT1Ds4FYa9hqKL1somb+8gc
AxzkFJ3Vk9enLz4HzTuRfobAuLoWM/m6SFYY116HIJeQ+WQD1Pj+p9FZQHgQRNYAEoyMTiT+Spx5h33PO1+Yy/4CgXT0zrO/smfeU7OgHiHLdmy0jfyW4+OZOgxYdKoH
GUnjBL5htQABe/EhEMqv8d50ZvHEhiMnsj/VPJPL7c5oTu2r/vCJvgdPbA8fSUY4SeFNNPBm8hnxlHp2G8L9kBTgJy3mjRf2JpH7e7WZFgDPpQevyP2E73PdeHSJPH00
8gednmzSVjd7og3+rYCNF2575JkGRk2bybi/3x/WdkKqa+371Ekbb0JWKOcKPmnqDH2RdZ2YNaP7I7sYFZEz4Y4czyK2EJDKB3EurdAe+gfzBODgyc9g1HPL+xrrJ+gn
XVUsIwV7m/crE/egF4j8fIUc5zAXPCFOpd5czvGFIhQcptjGmvEG4HiUMkc5PdkttnLrvRH2pLTHIoE9X+pwztvjC19jomqr26Uuv2Qsfr23+pVLi6r/cN5O+bS9us8D
4J1YnqzL1kKrSExJ4mUARVisWByskj5/vDXqZLmdpn8BVkDFYGzhcyg8e9L59u+JXNkeQfmSwgSzH5INy38r40lXQ+GRYKordTkDtdaestDPHH4YOFbqV+JTo0lCw+X/
pVd3zd04KWktD7F0hC+RxlpF+cL7/ySWffjyDtxMNjL5gMoayFR9FkKGPmN3CCPAIDa2VzVPeeT4uvgRmnvVsG9TgVgULaBxN2sT9E9Qutcp2Ok64vhAmCQ9ui345M6p
85yBiGiInO8MlBueHOsEXxMjnGxcF7FoD4asjxrz2Hq4UX57pNWuygLzbJtmqX/wymeomVncW3eySBocxl7an+o5Ku7pdapgY3tptCa4V5ulJshuvalJyhHArIhh5o9U
VYV0/JashMahGwOt7X+qhpiHv5CNW/CO9jShXsfqpe8iLJyOORNNu7SlbhXkwIL0fLa7BsW1A+XQPlLSMlhNj3b9xJPCOAW+D6WEW51ZJsFQDBsuKqqHS+Ih8UTGeg4K
7ORHPN3I4QnEDwvmPWk7fnILjpckxD9y2j3EhJVZVgR1OJQDFZBqba1hwAWtOwqH9cOT3nPi68WQpVuOiiHiFH1IKEo2SdJnyzr0362qFc6Oe+lWfnPt7LvTtWEql4Gm
RGaQh+QnKXYFHTDKJU/xNROqFJqt8v3zKv6b57MjWPwaQfTXr8Asd29RsYOC9NXaIRYemL1eYdpPRTv8BlXNJWYkmqYAhQ/hrupzHivVUvoGgyIc/DkbJJinnUgBuzjB
eoo5qe0z7B5PK3RvN/DS+k2s57Q86Wae8QfMbcO4Bz7KiCbRJr2HgYyrX3ljAm2InkPELMSQBI3KYVRngPExRizSthsSdYCUDp6Sue5InPEnP8w4VPJT8AuTH5BHu2c6
L6OYNbrfWCtP8QtppOVpvy5ikYiNpSLu1/ezzjFq4+vKiCbRJr2HgYyrX3ljAm2ILJNclFRv2hcb087cnjXEVFi7RZftaIQzxdKJ+LTfsT8Mt9N+4L5xLHYVPmSHgFqN
5BwJ5r0dhNW6F6o/grdZacqIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17uajDR93lq19jWzQidKggmtIjhPUODMVs/IQDPrkR3NXEpzg1lclRoRMSzwRYDFPi
vkYLX/miMK4iRpo4KSekV8qIJtEmvYeBjKtfeWMCbYj4RAb0fI4cA5c989xU/RtzVP3EylKFTJEwLexuvzYMbG/4PjLmHzWP5w0WYFJHI4xET2irJvzPNtET7T0SyIRP
i2Brb2P1bNYdqcrS0QfexHOQkSyvb3/+Ty8wZ34pJizd93Jg0pPUijZXofrfCAqhyogm0Sa9h4GMq195YwJtiHfhVAV2dy9zisaodInfmAw88E4FNlrLduaB0vosz+MP
2ztesKxOGtpVarBZXHKvN+fAfIvCERXvtTLZaT6qirYXZeYMJTp5dt1bR0AmYN1koY4ZFtMWUeI69RCmMkyCzQAekKIGLqxDIYQbcobAq0aFA7fbGcRKn/EOsH5QQNhg
00UGZTZVrfa66Wvj9adSTS536WTFDIpNI7Bv8oKTuB3KiCbRJr2HgYyrX3ljAm2IOgstFcV2Xp6gcZEZS3tvStTHu3LiE8P5N8Ennulhb5hgq1WQ1al/4sEkvWSq9JaG
ltLQX2u1qAfAEDjusK0alsqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOejCfNcbnQ8eC8VC3A/6mcJ8TkKwgTnqRX3r37atxNAwrM6MhjOyFIFTWHcb5pCtRqd
OWwR5mDkLZkDxdA26nHI7E9AHUqNPiKMXd6TmqYHnDF9NprB4chgHMmb1U5sOQsH7oFltv6q94Cj7iekm+tOV/kkpCLc2L9Zrq8SASdAHfvD8X61YgyvkbsBh++xi+mw
yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+8mchj7neTZr7LYVBpEOhzmSZXdRwN4saED/s81w/rdTIkX9yolj8/6R1j7soxeXk9cdTOXZQMBlvLrfa6IPB73
cgcuqXz8VKFxDjVJUfNjdg7c0lMQY6sPg3fnLl3PxCJyO94DM77/tTnxjBLslRoXd9Ev5tRQ9+bAb+QXcp3kj1yAOiDe2ivepRajyO12nmbKiCbRJr2HgYyrX3ljAm2I
UFcMrN2wuVtSYnoCCJUovAU3nbqNCtKkYgbZAxom+JQHiNkwb3IBmLCd3Z+7AYV/tRhNG+iS5uIUsw6feq7kFKY+elCft7zFIeZja7gl3NnXBJp0U5PYlRN43xU4ggSc
WKxYHKySPn+8NepkuZ2mfz1UOzxf8t+/3s9iPSEp38i6Zvj1DTAn3vpz8CVW14738wTg4MnPYNRzy/sa6yfoJ173QWpMSaXfNXMrI62u/V+FHOcwFzwhTqXeXM7xhSIU
8IhtFmjtApkwqUPdNxgWoLZy670R9qS0xyKBPV/qcM4gMw9oLcnVKL5HqPNKP/6748tCyOOTU9uQ5Mp3MuiSBuH95e7e3Y1jDiWM5+6Kfjiqa+371Ekbb0JWKOcKPmnq
JFa4ueuGSV2OAfl9KS7dkCfKV9yVcJH4AJOvnYBWGFoZSeMEvmG1AAF78SEQyq/xbx5neWCq13D22ZEf7iNP6TPvF7ovqAAEQnxiP/HGSD6XxX6C5/OG9EMOerGXgMbo
FOAnLeaNF/Ymkft7tZkWAFGt5DuZIndSeQWnKKUYBJUhtyfCIbvEqxtt3t1A+st4ia9fmNFgGjI/5LT99C91GrzA1+ENeB7rCIrRClnB3CDYjGA/HhfT94F0TDx7JJGI
jS+rCN1zw5BWEZY0X9AWCjORLQlRnVoFtwxPL0T1bCDhZxfgre0/qtM1NShGykI5LzGRnKo0BeEK5zuCsgHj0k2s57Q86Wae8QfMbcO4Bz6lEGXn5EpV9CcofEFEDkTv
CcBvhCSt5lzzPQLIGQ0EpsqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFz+JeP9p2tYw49WlVA2q1MJCqPZvSsJfn1fRBz/Evb+4r6gj/hPWpzJSMgZ2rvq5p1
yogm0Sa9h4GMq195YwJtiINxF05+fMMIhjTy+zEu7XvCBUmiRr5DUlYdsPB5EDX8yogm0Sa9h4GMq195YwJtiKpk1g1+NFLOKFDw3DyKaVTKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiFko4OuKoAYlK1ut68qYZFCGjgGTcIZ+07nkm2OMYKaAUNp1bqmHVvy30bZRA1z2/4Cjv0vYGEGhB3hfzRYrxHXKiCbRJr2HgYyrX3ljAm2I
shPhJeOCrw03Aj0EKt7hDi9iAkBTpDmeQbWg5YDq7gSwpb2MGxoBmnNsxN01YNcTpNfPngPwBpihgyYR12NLSedSoDfXyHuOg25YRxfbt9Jgq1WQ1al/4sEkvWSq9JaG
QyKgO+vP1DT5vgVhzOjJesqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOej4XS2Q1fnCtSLZ33wTlBaiMqIJtEmvYeBjKtfeWMCbYj4Lur34a7pZOjkr7y5BGsZ
Mkj5+YWUboWXRtQXctUCj09AHUqNPiKMXd6TmqYHnDFQDBsuKqqHS+Ih8UTGeg4KR7XJmO7os5yBZKBmGIwq73ILjpckxD9y2j3EhJVZVgQaEveNXwT9wybFp+VGzF4C
yogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+/qK476G9VDG4IodOsSwJNXVV9Am5N0VaDe4qxs+jMz8aegsTyDGFMzte7m7xEIQfL7ANa95qtwCohSIpMjnH1+
cgcuqXz8VKFxDjVJUfNjdp9eBDKziTdalok5g++VIDErlvR92lSBkiWuumWIQglwwCdj5rSXByAFXfdNDFRQpdcnimzwEO0GEmyJ6R+6ZJLKiCbRJr2HgYyrX3ljAm2I
UFcMrN2wuVtSYnoCCJUovM++2epGMnvfJPfayUfgZZGvb8pKIUMnc86CTcbkLt+zOYVsiatft+/31CXedmMNyKGhBBibOkZYDkL5Wc3evRQ2ZZaDXYXXaWDgGk1XVTzH
DaWsgj0D+ln2q91qcQ8yQDLhxmhYqgtFWuNBznYYskvy51hOGIZOnDR0STp9CELkcjveAzO+/7U58YwS7JUaF8qIJtEmvYeBjKtfeWMCbYg6ZwFlVR4ryg0wcPMsOHLB
ZRtxwm0A6N9usRQ82jApnbZy670R9qS0xyKBPV/qcM7a/7amaBLbDIE1iKuv+ATncPDIhS5lch4U3vcVL5HWWliDpS+0DPlIAX+Mxq/LEC2qa+371Ekbb0JWKOcKPmnq
izjoJo/rnkxgmsFC+wrUtceVkid6vefBIHJFFkHb98kZSeMEvmG1AAF78SEQyq/x2draDaO4SH0vlzWbDV/hNGhO7av+8Im+B09sDx9JRjjVe5AI0KMU8+nt02Irtz2P
FOAnLeaNF/Ymkft7tZkWANT6WCyE164HnGFIbJOulr8M28K55L888CVmb0+UBGteia9fmNFgGjI/5LT99C91Gk0RLf+jPdkbfLRQQmHl9J9EZpCH5CcpdgUdMMolT/E1
iBzAjpCf5bvKSPiAyUNRR7L9ql8pi252y7qRDKdV3sMNbCmqVmvaL93JZIVOvuDEQqo7c63zqZJXBkPdTIMt6URbntZbeVqMliJG2TRMHHz1Ds4FYa9hqKL1somb+8gc
TnwWdujCq0/qNb2Bb+jOjZ4hmRwdrBvDvUdeAs3k0BWqXU0HtT+eMVTl9oJBjZfXPvUdOfXibzV9DL88htA2RGscVRQbuNSp17eIXJI5C0+9rENtjWJHQ229BSfCYqYs
yogm0Sa9h4GMq195YwJtiINxF05+fMMIhjTy+zEu7XuyCHc6sjZy0aox60w6K2Y90iOE9Q4MxWz8hAM+uRHc1cRG1849/TeWFNleaMtqMMW+Rgtf+aIwriJGmjgpJ6RX
yogm0Sa9h4GMq195YwJtiCyTXJRUb9oXG9PO3J41xFRYu0WX7WiEM8XSifi037E/DLfTfuC+cSx2FT5kh4BajeQcCea9HYTVuheqP4K3WWnKiCbRJr2HgYyrX3ljAm2I
nkPELMSQBI3KYVRngPExRhhT2YYztKfQEfRreIOJt/InP8w4VPJT8AuTH5BHu2c6ewRCIRmd9fsmH288aAUGOi5ikYiNpSLu1/ezzjFq4+vKiCbRJr2HgYyrX3ljAm2I
ZOiBVPNUvrItI/ZJVIwN1fLuZQdyQscokSdiXTxlH74ahMa3HTKg2xxGkMFjQRGXI/XTKjHXCvcsIVzBR9ZWr8qIJtEmvYeBjKtfeWMCbYgAOKBfFkxQMNhXmiLkDRWR
TX90VAj5s2hN0DcK1cpi9HIHLql8/FShcQ41SVHzY3afXgQys4k3WpaJOYPvlSAxcO9FJ9UPSFHOhvdRrHl1wKaa3dULqwAjJq5GD1eonckr7qZX6//ardjeGERThQkG
cjveAzO+/7U58YwS7JUaF4Uc5zAXPCFOpd5czvGFIhQv3LDdW2d4LJrahPI2i/PxtnLrvRH2pLTHIoE9X+pwzrvQsT7fMjul1fBrefUO+M85bBHmYOQtmQPF0Dbqccjs
KbAWmvuvd8ilV1icDV9dy8BLGX1UQGGlSBs0L/OYhgkWMVak/JQci1J/FJS00RGjqTITzD8n0JwqVsYXapJMTqEbBGjpi76QB+2buigCleODcRdOfnzDCIY08vsxLu17
8ExU094L8HZFagC2u58nklMaEHlsnQsQyKZVFILUEq/+sKUxmHHllQCi+sYCz/W53gQg3m+nnSSytopLnlq8avusgKnLq+tC4WmAIYNPdvXodypqJjE7fF1O68p5RWZe
3s5Isej/I+MIwFhLo0puhWCrVZDVqX/iwSS9ZKr0loaj/2P8MZLiuBxBFcQVUdYuyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60+9VhXT8lqyExqEbA63tf6qG
n5RMGB2cEMCirr9o6qVWDpp1dNgiTqRyp45dhG2rPreX9/SnEbS0v3WJ84P0/ffww0pNaSbwTXJTrFhUYnn4H1isWByskj5/vDXqZLmdpn+5XQhzfFpT/tJ0IV7hN54l
zRG59FbluhV8VHm3QS5jOvME4ODJz2DUc8v7Gusn6CdMKn3qo65DYlNbf2a/rm6QM+8Xui+oAARCfGI/8cZIPpfFfoLn84b0Qw56sZeAxugU4Cct5o0X9iaR+3u1mRYA
b0J+UEEll2joIPVpqjBa9+wu5xKqB2VNEsxw7AOyEwmqXU0HtT+eMVTl9oJBjZfXHchFmgaIHR7YQJZ/DSR5nFMOV4zAEkzbjrg3UC4JbS8sG9ai4+jEsajDHj6zYD8v
l3IE055EmYSwZKuGIhmqYet48B4+Bk09Fg9hYF35DqJG80tRaBVFIPItqqaQw6EYyogm0Sa9h4GMq195YwJtiMRSIllXv+GPmmydc4i9WkbKiCbRJr2HgYyrX3ljAm2I
T0AdSo0+Ioxd3pOapgecMRKxAH3sNjMnNXoJcwF2Iu4wzRQ/IEAu6lPvglUzIp4s2xKVbWglVvs/Qum5AlqAts/jmypnhhqUpF2dZQyduprKiCbRJr2HgYyrX3ljAm2I
I/IDSjaiRHEemtQ1TLV1v72sQ22NYkdDbb0FJ8Jipiz7GF3hkVzKZAoM5pJGg1HvTACawx5ilbhhZ8ahmwP9acqIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0i
htAcn4WHa060ztPU1McMui5ikYiNpSLu1/ezzjFq4+uPGV0C0HpjXL5OOg21PLA/yogm0Sa9h4GMq195YwJtiDRYlTE78nku/iN2dKkUNF+blAZW9cvhIEl5Jmy0Fh0F
Qt740ybFOyn1xxQWFfZN1X4RP+VDy1f8YAYz9empzSHcO+XZTBazxQZG4eZ2cxsTQ0vekNgI13b+cHi6w8qIVVQhKtFhnQtcwZLZFC4Z0mQgNrZXNU955Pi6+BGae9Ww
x5jZ8kFvTV4eNUYf1pBM4IJ25f5Bw+Lu1bVQPXIVI8TE+ntwyPx3mOepNIb4jB5oAxzkFJ3Vk9enLz4HzTuRfrSQmYx7t7RK/Jmdt0JtAwM7aRiHyyAhBTD0bKMRoFJ2
dXxXtVCSZDC9p2uiSLlJA8pnqJlZ3Ft3skgaHMZe2p8bX+469DnS50B8CPdwzLqicF/B5flQTNbVkcJhs1EXQ4EVxi5VlAlYBlRkZqhd/moDHOQUndWT16cvPgfNO5F+
sEsHb3NfTLOc/ATEYaPEaiM+VMlz5oTs9LOu6rO0XGazST9yH9RxGS5V41wty/qqz6UHr8j9hO9z3Xh0iTx9NKS43pZoj1I6yf1u16Pc3mo1OWIIES5dTOECIF57l+fS
Kr99Q8VeSDlq93OBLsqQY8+lB6/I/YTvc914dIk8fTTs2WevfC8Mit4y2CG3HwQlIz5UyXPmhOz0s67qs7RcZpVMjnrK2jxh5h4ejAWtqznb4wtfY6Jqq9ulLr9kLH69
POjYOj9BZWrQ/LXI6SCUc+gvC3R2GLp1uSzj7iV6A3RBTbqaqHVnlIam61jD2CTyIDa2VzVPeeT4uvgRmnvVsK+atF+neevNgOIxZrPKOfsjs/aWPJPXObJoYLvMzBmL
G+m4Gy88NW9RfmZJuqa69iIsnI45E027tKVuFeTAgvR8trsGxbUD5dA+UtIyWE2PitkrTRS5xgaWcgkB2y/MN1RJ94ro9Mth/k54AftDQPUAtjW3m2rtRD88YdozTcLJ
GUnjBL5htQABe/EhEMqv8XYA4xSIHqQE2ON1iJMin0zTw1WNBrl5zMgMVfnZeYX/ALY1t5tq7UQ/PGHaM03CyRlJ4wS+YbUAAXvxIRDKr/FRWOJAnqZl+Z4y3n+LZS6c
6SZ95F+hMhjivkInpIpilSrxH376J1gkYG5kJNmHkD7zBODgyc9g1HPL+xrrJ+gnYrbAI2D9pks7dh2ykgFAAEu3Vri+liEoGSD9vARQ7rJqrhay4gq7hsSMb6IB8RZR
3Dvl2UwWs8UGRuHmdnMbE0NL3pDYCNd2/nB4usPKiFVngyeLfTVohu9EAzu70I58IDMPaC3J1Si+R6jzSj/+u9rOGyZsI1Gj823nKtdPCvZa43zOUxFI0q+5a36QZKCw
ZpybsZrXNKq40Ho4H121fHy2uwbFtQPl0D5S0jJYTY/02n0BS1Jh7S0nSamh15e4Om7nmn5VkvPfMjlGZ9uI3ufAfIvCERXvtTLZaT6qirbT6E5Nv8/9H8yn5zTB5EUw
F8Mtad9FAmBDWvD2JdTR/xV5ECxGQ9AkfELIrWkEpWUMYDxYyaRBv2n5LlYuegIBzuN02sK00v3yW8ipwPhfOpkOzFxaDfR36N6xd69vdoH8wd6Y7a9cEapX0K96FFHW
8wTg4MnPYNRzy/sa6yfoJ/+eYzXyacrayGcaw/mwa/8YXqG/vpA5y+HGZ3qsCyJp5KSeXsPzmGalKqP3dNvygVWenTDCmra84zjwxtBf2iEfuqyez7d2uhs6v7M6pAhb
KvxET0tLVGCXf0deTTFJ99SQfy9eaSUrRdRyOCDS747Q9oc7z1AzoG6bh9Xb1B9uC+S4+hoxqo7450VTXWtn1tBkQx5CDkt36mikPH9a5bkVF7wyx9on/eWFQRwzqlQJ
wqPw5CJLYUWWRKkmzXhu74JokqBXtK1QXL8VCQQNq7s5hWyJq1+37/fUJd52Yw3IEoRrYBzZA38qvvQmva6toVoIY+cp2x6UrTrh7ixoO3uBI0kJNmuGrF3D8f0nWenh
1JB/L15pJStF1HI4INLvjiQcjbgRGhZzk3Da4HbAFZ7Ay25oL6A0XN8jo69Wgd28KBMzTuycx7hMPkQ0nE6mjjJ0bH7CWlSxAa1pQ9kHic4UhEZNHV36u6It8whLTE4C
GGSVeawfzRnStgzb+Vu+shi2XzBbf5kJ4G7Maywg1S9luUGxSFMWPXZBYqawdfPOsKUlBo5sx1CAEasgv/DI63n0mkasGvkT+BYV2HxD2Ka2MDkmfcxoydmbjXXANtGj
0+hOTb/P/R/Mp+c0weRFMNmTsuBcR8xpGHyCuGFdMeA7vpLQU/Vj2Y5EIY3fS3gXmnV02CJOpHKnjl2Ebas+t/QvUWpWPkJl3BnmoXrrR++YgxudUOVV5rpbqIpCHayv
eyO8Yj0bLz9Xi4pgx3Q6CKo85yIBuUvhcQCxY3yKk/pkjb7owkbC60XvVJHOWzyUfcm2hG+IOPXPFN/6VeGMmSft8njzoLZfJkjVEA3GUoodDzvCjNT77i2NpjkAPOm8
Zm1d3MC3JOjUnf8H5vX+seu9iSp6hfStMsJxhHyV3tWQl7R1G73J1Kx0A556GbKOT0oX2oSDfsmBg3GoU0Zq08oi8JXzLdmIr5+bIa9fc9PoxLK6MGnMhqf+v5PRiZ3z
gKY3HOKtNh3t9dyzixdUhFgF9GkqvI3T532KH4N1qB0MdpCgTqnYMqhioRijnX9OWTA8N86wIl2HZajD3Qahb/2LOoTQakhdSery41MgGwSgl3lSRxk3S6Re5FSFEU7M
SgEQuSBNhFMpCWNGJR8CheKvwfDvNMfswJomrSPIH4alcoewlXRiquRtcz+h3yI63mR7bwl6s3I5XhA0E5TXqUWPGTW1qDVZ3fUtGbxb9m/K77RB6IEtqVOQ2ENBHstx
V0qtsc0oR7X06bTRgur/mf6lDkKM06uwSI0qPfh+/4y9ZFQqpWEWGQtO/+ZeSBROMiMvU5T8ts7YHaviRNyHV6y7AieKG2XhjDpp8/u2lNd7se/oiXmQ6yyMkp/1c5yn
a45AQE+CvRbtELf1zPnponZjGx3TFv7UZIuRtx6ZN/MtKa2m2zfMwXWoCkAXTqs9zc6q9uiwWQAz+ylDVCtFslWmCXoiz2mSnKQrd4IEuqLe9z1qrEwZ4WloQ1nK4n2A
/yvC+eLUVgi99hR0h8Twv+hA1A7NfA8K4wOiKxijzEAujnbpEEqNMe89IsafrMdUa+5DLCzSOXS2+IrNyQz5nFtrn1v+hXO4NVidVts741qi/vLAQGJw3mABeXRVY7IS
aG/XZXv73RO1DZUpu3iNb3Ne023xSfiU+e0y7JbucitQ4UnBkDIrATBm7se0jqV89JovoGR5GXaN31fADczhj2EW8yNkAhhGNQ/qptpaKgkg/M+RkNBRiovharMAYzTi
XO7hHnk/duC2aVOtdfWehre9nC5YzLcsGyNxdRtOawotKa2m2zfMwXWoCkAXTqs9zc6q9uiwWQAz+ylDVCtFsnTvWBTNw2jHjwFN27U2d39Q4UnBkDIrATBm7se0jqV8
HE6t1dTGrSYngr6zsHvZi3GDPKc+UuwwsWOcfFAt8VGolGVKtK/6ceVvqkGCMmBVSnjxu016IOLucmLeLDWKef5Y0IrBpttDMmPH6IkfPmi+BoKscjiS7rnVa7X4PYIq
Wjlq1WqUffyINlrIa1jTSmTJpIwpxkycGRJsy7JdEuZAnLHmwpJ+Y4kojhtHL3GVnWN17tzWfU/U2AIe1shYUbOfjobjlRzLG0dh0w4iq9jijJr3D21a9bgoc/xko+/y
8MP2BP6E8PiXN6yA11NutuEn8a2nOmEQQUvLv/ScFn1KITSbTYJw1RHvwvS2sFVEPdpfriBenMSWK1fGhYYrzFLHolebDXbIldxnP5shBNWUikjfESqnwO8T2wHXdLr8
UvdYUCmDFMYqebDvjIStfKiUZUq0r/px5W+qQYIyYFVKePG7TXog4u5yYt4sNYp58aueeDpm6fRHb1mn2YrYv4ZOjDhxYt7DFVkUIClERxWLJ2V2PvCiEGEO+KqrUptQ
Bahb5reYvqXahs3up4fh2xCJLOS+HkbD+vejgUAUYcEjqFdNS+/ooGsJ25OPs02GCovutB0rGq2+5CgXUXGBi3SbgQQb2ZUnXt1YTk4A5n8sGonh/WlzTvAzRlMQ6Jqu
ffeGBVnUEGguqlbZlj3MFxdzdryIUDjmPnB2blSe6/XGA/02EN5Nf9iZ1874BMG/gKY3HOKtNh3t9dyzixdUhFgF9GkqvI3T532KH4N1qB0MdpCgTqnYMqhioRijnX9O
wt/9NBX3l9yZ4bAwjTgZ438j8p+UyDkmlhSueoDNYJiVfffLhyPV/314E4xbprSS/nWG9uyZjBYhwnJQHXEyFg1CVL/Ux3Ipd2eNqr1Et4MjPlTJc+aE7PSzruqztFxm
1y6lXg0iQWVwxwpaJIn8IUAddOLvG0Wb2DHvruknYfS4qmkSA7rhClXHUpttuJ/p6uk+2X78nvZKLfTL9nZfv1i80OU97Vjzi/9DEns+FmC4qmkSA7rhClXHUpttuJ/p
ZUPby8O+y67ytsTMb9IHwVAdFwwTh7xX+HNtnvWqcq4jPlTJc+aE7PSzruqztFxmoFomZl3bNDWm8zPHadYUtFAvmKEH51EDlNiq1GNr+ZMjPlTJc+aE7PSzruqztFxm
hFHhq9In6J6Lg6wFF4yjoOSrXrxny/2AeIMBc4EpUGheL0PAJfkR+fgEqaLZf0GOZkUJBRJnpdN8sKg7l32D3Jp8W11fOveDKlurisfKtwEZ+Ku8h3OyghV3xCrt1/bt
U2Mk3q1wdLLtY2HEpSfYInZMpW8YYhYIrc+Fv6LqEDTDAVEi4t0nOrEe04ujexFnIz5UyXPmhOz0s67qs7RcZrHa+o9IVPcrQ1AjBb237HxFFYM0p3YH0lZ7bpzWjUU7
S22E4gg7fIlH6gNoFoJ0Mjw+0gMcegD4w8Tp3atmH0jV6AD25bUCmhB6EqqdUzYt5RZk8e0LT7KPY07C6ruWogxho2El/5iYVGXTBT8GY9a5jXdUKDY/uwTCMgUweq+M
CHI786yrDnnTnPYQoT+dzkDWVHY12L3aOi/sS0V2MFhKARC5IE2EUykJY0YlHwKFj3ii/dj8aRWPmYpM2IRdnwhyO/Osqw5505z2EKE/nc43PEn7mVkNmoSTGqIWfCS5
SgEQuSBNhFMpCWNGJR8ChawyzAOh+UKBrTQSgRtFHsMIcjvzrKsOedOc9hChP53O3ZxRf6QF3YOhXQCMrdR0veiKupfWzAyMYMvt28VMBdvIyS2M9Yp2YfSPs3zSsS3+
uKppEgO64QpVx1Kbbbif6ZCJ5JE+YPF02xH1LbNuUCp2OMsbdUIHwisWTrl8dzQRkInkkT5g8XTbEfUts25QKoYYTDKLLYzITi3l1kDCq5G/F7SPlj00QfEG9vyk/p0+
PQtD8NafwSyWaYXljkc3sgdtEqt3chqGi1MLMP7IpZq7DmJnt4cVHEdiFI6rCP/wvxe0j5Y9NEHxBvb8pP6dPlfQkvHnA6HcpmkbXHR8ZJ/+8jAyvd+6sBabQTFouHkf
CKC/tTfJC1lxo2A5U71LfEI2A1R78JLar24ix97M0EFxiKr6uFRgofFd2ysmM56VFXnih4BybSSj5IapNULV7JCXtHUbvcnUrHQDnnoZso62XQo7cC793zCz5ylHnM1r
T6Z/ZeQMOGgudhSLEaTWClPPSxBcfcxVu1XdxnPQeUoaP44p9GQ/FJ++OsbLOVrAZI2+6MJGwutF71SRzls8lBQfg50JGiSFvm8Yyg7PO3KVmEA/6lu1E3JDvTp7QAa4
wedYTg+t5Z83M+ce19jArqp6VdbxhiY/zVXZmD5nDVdEXIQX2dM1SfHh6iR4XR5pyu+0QeiBLalTkNhDQR7LcVMxyhJSAwpj8KjUw2kimH+x2vqPSFT3K0NQIwW9t+x8
/Ys6hNBqSF1J6vLjUyAbBKCXeVJHGTdLpF7kVIURTszcVf3v3/fqeW9UYgJGjcCxjFUYIbTrtvL9h+HTQcHFhAA8zi0SMruJiw3m4wuAjfyPNslFyfvnJFkk9DW2uFwY
0UuhlA3PO/Njca/ahiW5FYo3ZWm8yuDEYCDdNN+a+wVrvmfC0bStZKXmrVGhpYpYsA4T13tEiXEXaBjXgDII35pTgc8UFg7qHX2sgr8W3I/B51hOD63lnzcz5x7X2MCu
qnpV1vGGJj/NVdmYPmcNVxdt12PBKYjBrtdScumn+ZtQ4UnBkDIrATBm7se0jqV8eednrdt/LyamiZGxjLCYBYrPZZgcPpe+C+R9l6GSL374n2H4qi8YEwJhBr8yPk73
bBNJSZl8taEyHim9cLp6pYuZrFOw3+zcQHHNuaOH+/U5Cf7PbuxpOx/n+8EYnKzGZzHu7ulUu4VuPROQlM02HdBzUDW6wAzFbGRMhw+I8wY57qRqmhxNdfnLS+SNexBy
NgddiAv7JwO6FUCNzYfPbltrn1v+hXO4NVidVts741qi/vLAQGJw3mABeXRVY7ISqwohZxqObeI3y0/1/wQLMQP9bEmm7ptGufiEOwjFk0oKrLaBMBn/wRKBSaGXawA+
MiMvU5T8ts7YHaviRNyHV1daHuRLua/3tZffJYtePQWJ20Yvj+O2xBF2S+9TqBQ3Oz4VyjAcg9Zlj+cwFwFDXjCSH5PmcPvqeOyrDztKC3Mn7fJ486C2XyZI1RANxlKK
HQ87wozU++4tjaY5ADzpvAyA00MqQ006vUFoPtyL69+Pku3lBRd92YBUx9asJzV0iydldj7wohBhDviqq1KbUPL/wEZmxqfX2LdAcv6A7r2b2BNh55TQk+b8gwIF7NFp
9JovoGR5GXaN31fADczhj4OfXTgTf7m1EhNPxyIsy675kziYotNPnbcFj30BaAyP2suyFT0OyDthqmJaAr2uKXuVG7DYi9PlXFAGnuHqrUC1a0cJACAyhCvjaw8ohykW
yu+0QeiBLalTkNhDQR7LccqBgCYD6db4KMRp+bCcZyBZKqT0E1yLFpnfLp7vBuOrHFr5Vvgg+hOT4oLzq8E1b8Ac06GU1hj9cvxxL0cXVIpvC1mPnNiEQHbdY623qZlV
I/jooot0bvq+VVQM49CuIKgPeRSiiiBSLrNM6L/oJvYz6Wr3Q4tCBAJOX3Wk3oqTIhHc/mngAQfoYgfaZyqwzZvYE2HnlNCT5vyDAgXs0Wn0mi+gZHkZdo3fV8ANzOGP
g59dOBN/ubUSE0/HIizLrnux7+iJeZDrLIySn/VznKdrjkBAT4K9Fu0Qt/XM+emiax6dS6LfqcbMOMa0SkCNaZNN33Oj2BdpzaKaV9WGQv18hz4sViIAFjhlAXnPznmY
s6sj6OukgO7Udz4qPWU5mcBHGkdCpBEVFc+Y9V217TyQl7R1G73J1Kx0A556GbKOGAMg1jSSDJ7DJnpkMrq0i2PimyZJR/F9W9o3plNNX5Hi4Dv7dNKIYpXGEPNIkCuu
ujKq7Lb5ixh5cG+KtsY2C/WtXwa4b3ufmWpW0JFMQ6SCV6Ria1NWWPreue+ET2ktowBBSbOur9WBNIlumYw4+TtMTIqJ2MadmFBnOR+Q51eAUqHQTa7h21GH6ln5Ld7e
oDkxaqYLi+aiOQ+yH8PsdA7f6diZ6LcPrbzrI1dj4T2+JG6zzXZift5o3lAtSV8xkJe0dRu9ydSsdAOeehmyjqgU/nKyLn6ggY/ctkyRuVn4n2H4qi8YEwJhBr8yPk73
26jbKj/5pfy2wm+asRE+AfkhF52BYwckfQ5GyWbYOr1rjkBAT4K9Fu0Qt/XM+emiggSGh2MvvlUW5lmo/VfwtL4kbrPNdmJ+3mjeUC1JXzEyIy9TlPy2ztgdq+JE3IdX
7xNsfSnawPp0418jdqIPWJ15LTrKQdfasgkZEhMc2QG3ocA33Gpb+4w1/jx/e2VACYw6RehikSpWMnUeb5/v4H3+iWyfCJwL2pzl7Io0ges4XaLbxzNx5fD3BpaHiHO1
vg6o+jP2Nx2UMAkhgwXeaK4WVpCiBDWk3zRHo1U5q6aU8U2PflUgLXqfj2Aa9baCtbh3hpeNKr6X4fMOQW9GPe8TbH0p2sD6dONfI3aiD1ih/mbFMywvnV+gR93qCJpb
MO8Vs7f4vqClkNnkiO+dLwmMOkXoYpEqVjJ1Hm+f7+A7TEyKidjGnZhQZzkfkOdXy00CmsMoVk6tKs0GddplG65XUO9BHJ5kC2kfHzI+VlmZqKITP1UFaaWNr7TMlZjt
sL+l5ixmlP3W5K+q2vbiZ/U1vdtRhVL8t2jhUaXE3/Zgve8ymNkD947ZoOaO/rwF28Z2GCP+3syRRzBN1WHAE83OqvbosFkAM/spQ1QrRbLzxrk125SroEe7rVHptfM9
3vc9aqxMGeFpaENZyuJ9gEEZNVF2zpVXFHcYzkKIaFrhNbuCNdvw/ygK8P5hdFIZa45AQE+CvRbtELf1zPnpopJYF/k5E/ww/GMZT3EaqUZjHVakkbtYP8iLpG2slYx4
IjE1GaB+QnvN5t/w7sK8yvxe3ys/Z7A0Akzc0zSOQD/FXsZZIzYcWW8jfy674uEWwedYTg+t5Z83M+ce19jArlL1bVEYSLCZ0J/fAabV6Bxba59b/oVzuDVYnVbbO+Na
hb7NBUMJAj5WnkvUVcUuPcqJ3B3DNwhGCDC0chF2XfxzXtNt8Un4lPntMuyW7nIrm9gTYeeU0JPm/IMCBezRaRiQioVVj6lgLGOCqVcFvahhFvMjZAIYRjUP6qbaWioJ
1QnqTEnpyXPrwpfLsoyEZ5/4aR9iIhqUzLBjfJYT7e+gR0A31vcJw2Q2KM8LRSdkHQ87wozU++4tjaY5ADzpvCgrhw4l4mfPi109dIgmxfMxYmf9TfvieZq4i1+4laBe
+/PFJGZZeY4WkkqcDzxHwNJMZ45uzt8r0f/MToicFDlaZJU0hHuB0SDxDxMB4K/7HmcEzAtP6wSVwuUCrOrzcE0CfvgamVFeeL9aDnfzJYwgmc706pqpGQo421FyR4ow
rSvchAhyyW4vArGqI+YlD721jSWOnkx+HKg0SkmdrkClGesFthbxzBs2DsF7/hkXxOicu+hDEiIEz8YgH2KGt50WOeb8VcnGpYEpxsx/eXdShpIHg/AIpZ7VhUJ7hkw3
u+a1SkC9jCo6yUmSpTNeIjklZvoZ733LOevuGEBLqZDe2DfolkiNM3wPtVD1H9WyJiRUGOCDC49p8OJuW965+J9W8M11b7bOFK4KletK+lZPij7JwWM0tqL57l8VlYPP
t7PhCJJPp+5ucGgQPLSVKC6YWEfM2QquS6/bweFU+ZrH9O/Je6x+Vp/Pkztc/Zy+yAmBtRdnR6sw+lSd2UIW/VY6Ik8kmnTTIOexIVqXAG8VUO2lNZ59BMdS+Y009aBG
Wazflag//GrTi+1JwdCAVkmUgCxpWYPbbZs+0fwbUt2wV3jHo5iQlT2fx+ukkoURrhZWkKIENaTfNEejVTmrphiN8DVUgmjhxj3kU/2jGe7+q6sHqdkOWMq2mOO6rFmR
SFvrOJkeHsrE3695mC82BvdYLhW7PE65oVxPMtO3wGeTKM1u+2Wg4xOxaWGRQL5KyoVS8/otjssCSEzyEjBKN6EWBshvp6LsGW+4Tp9zwAXuOFfVyQIwdFkKir0gRyJ8
vMIslQ4UvLVW78fmANDoUBqlLUXAIeWKwKwtePFcjWzzHfMEH5w4+ipclzy56ZxFwGvCxtUR+SumCx4VdOL+Mv6rqwep2Q5YyraY47qsWZFIW+s4mR4eysTfr3mYLzYG
qXghEQ7eaItwNKIaFBqiwLmOc/1Ih1KsLB75jq5XqUSn7mPN3n3vbxrh9R6TyuUQzGAs+hT48tjNMh99d1Svuyt4yzJRwMwbtPp+vPYF5BG3s+EIkk+n7m5waBA8tJUo
KeMfeJ/QP52UlB2f6yH5Ak+KPsnBYzS2ovnuXxWVg88K1N0vzSteUeQmGHCCp1cjWZM4SJDT2+G59mTYe3BtDz0FmkA9ayQe0VftGiKztVz7WZY+Je3TftHjcweMBxeO
+/1aquhJmcR11K30FjHizUmV3UcDeLGhA/7PNcP63UxGg0Xugm18crjVFne+LKExUxoQeWydCxDIplUUgtQSr94ER6ENG7m0FDD1bgBFTDrcD8dBQBgcZjBz164qcx/8
9vlM2Ki0cwaZftSjBWxx28qIJtEmvYeBjKtfeWMCbYjnlc0/TnYDMr52ti5vXatNpQIDdhXuuIMkKx6nnKL3nsqIJtEmvYeBjKtfeWMCbYgSRqiVp9bf6hq6IpjBQBhW
M3RtMrLu9G94daKazCv8YkEmaUhTtqNXgLqditg2MJeHuxxrwFamaVBSRfmiZzyiIbwT7+LM6ANm0JxPpJjbxMqIJtEmvYeBjKtfeWMCbYh0QylWTT+JUsH9dzyAo74D
fX9Es0IIcMeEUy4m7v+KRmRJJY4rk7InR/dwo4V7KRCHTGN0jDrQ9Q2H0Bi4jnxfyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj2uzAflGXdSR4nP5/retPv
lYplnaKjfaH7xzeC5ZPlJLGR25uA4DJ+DIjFkLkytMXX5VWb7EIdIAQ9p1+igM0Zx+1Rtl0N6vcROnBIrbvLPgQkgHhgJpwSdmaWWp3h246BGsicGBkPX0c32PkFnOej
bRNG8BFa27XntGmIAMcpct87eGsX6gYkvacBj9HvdZFQSFOgCsOCVwMnd6Mw+WmbD8Lt/ykt2+ata7FGEh1AbVAU4bEI5ktLq/lx1MzGeZOeQ8QsxJAEjcphVGeA8TFG
0dRUcW1kBN0QP6r9AXUH+JcwINzbk6I3U+MBpTF9w5sfuFDfIF2pOXQjcM/PNiU8sA4T13tEiXEXaBjXgDII3xbN6GLy6nFuAA9pWFXyf96DcRdOfnzDCIY08vsxLu17
r3BHxdEdPsnrYsA3HT2E8Och+xtdBRQtczVnFSAzdJPZuc93f8fglnPvvlwNK3mppDAixgPdhmk/Wm6tR3wtrARbNxbxf+z96yrCQzSamr/TIZGc9kTWzrYMDyDvnYgc
80s1u2OqHYTm0Fd/2Mp/6ALEL1e0VhbABdRz/ahuEzEqdq4cL52YJJXsGrzl2U9l3FX979/36nlvVGICRo3AsTUOwlGmGm4su+hcsCjUHazeBEehDRu5tBQw9W4ARUw6
3A/HQUAYHGYwc9euKnMf/C98GAo+SX8g9NuD4UKl/TzSQ43EBgKroxSYDs3ORJtMCrOzsfJW+fzZF8vlU3DWkd2cUX+kBd2DoV0AjK3UdL3KiCbRJr2HgYyrX3ljAm2I
bcx9A3euJafUPZh7l1vZhQ3N7lracVCnElWQT0pZJPTKiCbRJr2HgYyrX3ljAm2ImvtDOyt68qD6Y6SaxhVLYfPCSoSRKXjsEcS7o+InP0XKiCbRJr2HgYyrX3ljAm2I
dEMpVk0/iVLB/Xc8gKO+A5fXvBRS3lpfMexoqRZkiUjKiCbRJr2HgYyrX3ljAm2I3HfMce1baEkNXi1VMe4CxilA8KMxvnE/m04N14URnbhyO94DM77/tTnxjBLslRoX
QMmqsJAIM6uAKSZME0akDD+GaeXuDp5zPy8CFEmAMYEkVri564ZJXY4B+X0pLt2Q9Q7OBWGvYaii9bKJm/vIHDxYJQPz6RhUoXOVij+5WMDKiCbRJr2HgYyrX3ljAm2I
gRrInBgZD19HN9j5BZzno/aPXX832cy3L6chrKxFaKv7/rAclfuiqXuFWRIMN+x83kENLmSi/T//RctpfHrjxsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
nkPELMSQBI3KYVRngPExRj9u+1umbiDECcOWQCCuA8WXMCDc25OiN1PjAaUxfcObfvKjfc9lnGu+e90XkEwvwdSLMvYG46NnqBdqbcM2zyk3pcLnZ9blzPtvrakIynYD
g3EXTn58wwiGNPL7MS7te8iDUGhKFkp79ZDQ0AysnhrnIfsbXQUULXM1ZxUgM3STeNFT2P/SNF2QbwEqN5AtMeEiqi3FWv+mDG/HBYRAWcejcOUA4yoCLOZPRMdCiJfz
Jx7JHwfULrDpdqo6GODMdvNLNbtjqh2E5tBXf9jKf+gKOp7bs8Jy9SE2sLt5cE6Gcb31qIW9u6RLwqfJbPatvHuVG7DYi9PlXFAGnuHqrUAOCeVZheSei+2f7ULUrpV5
ksVCEwYQqdTtxoDIQbz5HdwPx0FAGBxmMHPXripzH/zGu55rrzF3vSDx3C2DlDbXpMdkvg4aePZ6Z0eyzw0cIs6wUuaA62ahqzL93RruLHyoO47DyXYZ/rK/4lGYa3iG
Ms6Yp83sbEijSPVFltsRMG3MfQN3riWn1D2Ye5db2YWFoMtrUWJ9rZ6leRSSxBmt6aDgpvP4NbNauVvt6Dfx6pr7QzsrevKg+mOkmsYVS2Es/5+QaTWo5sL8wdEAA7Fb
Rdy5PvRglrwdSL+aTHC2TXRDKVZNP4lSwf13PICjvgNrT2aLYrE8o94M8Rpyn9MADt/p2Jnotw+tvOsjV2PhPXGopaQ4sec07vvne7kteS+gb5NCX0h2/ImG4tzBlm2A
5c3YPwXRvIsngCSOjW8VY/a7MB+UZd1JHic/n+t60++0Jt9pHP5OKwbdkUDzEkXVyogm0Sa9h4GMq195YwJtiM7NdkBE5clprS7g6VxPhU+Ps0lPd7N74dCSYVTNAkvT
i2Brb2P1bNYdqcrS0QfexH1IKEo2SdJnyzr0362qFc7MLIHCa5GYHpBy+T6fqyOvyogm0Sa9h4GMq195YwJtiBTgJy3mjRf2JpH7e7WZFgCBJ0oShq4ZEuIe0pO0XA6h
yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUbpcVYkOJUkr977gqlum6i6LmKRiI2lIu7X97POMWrj6wEk6acOqOIjL07EDG5KKKlzvqC1TQSMcStr1RELn61Q
2wcJG0V1nmsEC6bN4/QREYNxF05+fMMIhjTy+zEu7Xv3Vce+AIwqMZD9ad9ILfUkyhv2DAx6htG2rwiEmWl+ZSaN9KqRKMAV+2HiwOPLtP1WOiJPJJp00yDnsSFalwBv
AxWfTmo0VNdz/UEl+7m6PPeejjX5LVfeAaZ/Z40rzhWSNw09cGng8UC0zuarcnzVgKY3HOKtNh3t9dyzixdUhEmV3UcDeLGhA/7PNcP63UwR7Q8A4c+Mw5VXgIj1T88O
7VzB24ecJznOUmjC3bBU2pWyZnYRh4YEStkzE2V7Yu0rT0IBoL4Z0+hOhwgDG/l47XuywOt9WXchxxMQsYRjGYlboF4Jz/nIsHVOegbO8h3nlc0/TnYDMr52ti5vXatN
LphYR8zZCq5Lr9vB4VT5mgfyMVjlEIvJecvAy07ZO4USRqiVp9bf6hq6IpjBQBhWw7/w+EoArVCloHhVvf3ZTYU5cdRuF9j/DbP54eKnvCcix/tmAPiFZNwedTdnsJDv
g9iy0PJ9BibEsGkeRJrRjffWrL5U/CNEWpMnrPZodjEV0mRPfb2LsI6eEzUpjEqh7VzB24ecJznOUmjC3bBU2gqOyhoKxJaGCt4myMNaNZLcd8xx7VtoSQ1eLVUx7gLG
q/B0cG0o8QqGrpx8QT/Xa1xvx6iadwKbt944LUMspXFAyaqwkAgzq4ApJkwTRqQMZXdqqSS5R3O7muBF2L+sg65ehsxIxa06CYZd1n8TBffOzXZAROXJaa0u4OlcT4VP
SiGdAIboKY9SXPzUKSG4WyJdTb2+e5138jetHbtSKOi+f7/TWd+gtZE5vwDxIiGTHcskiWWRcAwAB8VxdE6JLNO9UcovqogNB4XboNXjZzYe07czZ2duKjmUJjU4wmLj
sFd4x6OYkJU9n8frpJKFEQ7f6diZ6LcPrbzrI1dj4T1ugT+Y+erPn+0N/PpJCLuHITNdVUc5/0T+V9SeqHZ2j8qIJtEmvYeBjKtfeWMCbYgBJOmnDqjiIy9OxAxuSiip
pVq5uKrvX43QT+Ohi0JJ52C1WuHTTa8CRIs1N9xZRxWDcRdOfnzDCIY08vsxLu17yAqhGjr2plpnm7Id+8x+2tb+4DIDIei485raQvpUrAEmjfSqkSjAFfth4sDjy7T9
ZVNzt8QXph95uqya53yDmTRoQAgq4UfbWtCek7GAQFXTIZGc9kTWzrYMDyDvnYgc5XKuS7fCBHzQuCryvzt+pIiTzaeBQzdz2bF8pd5cNDJJld1HA3ixoQP+zzXD+t1M
PvUdOfXibzV9DL88htA2RMqIJtEmvYeBjKtfeWMCbYjeBEehDRu5tBQw9W4ARUw6zV7S7XwwEc8JlT9ny4w6i8nw+AIvNgL9Wp2Cl1L1ay/KiCbRJr2HgYyrX3ljAm2I
dU0Pjvjar3qxxOFipGFJW8qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IeYaRd5UJvhATJRqqCeer0zjPVMipVwdAUhgVCzlw4rm3AnAmr1DpIWr/eE63BE6l
nB/u/RPRJ3uzKuzUmfikf2xKVlVH4eDW1Ah1R/vCYO6xZfSJ+4r+jcaub6tTgUpXOyqVspvb9GS6Jyg5BE8qERxCwltjONpvlYBwIld9R469J/9vILY/7JxedG1gBtpm
WKIz9Q9vwx4R442Tc3bJr+Hk2LrhAANW8003om5Ytt+efXonmki7Lldk05oArVQanRu+6k9KS/9uQT10PQ6gcnyx2tTnFV7s2W32U4+lL7O2EA7BluYntf3eC3RHH3pC
X6X/bony1E84461VK2ul9hyDQP/M2RtjNlvZmbo5mHEHkODPDT5wKMzJe/8TUH2mqKmknd5E55lpEDp9sa1AZSM2t7syVTaOjdI9zJQADO0671rsJLeW8Tn8sqMfIBRO
GqUtRcAh5YrArC148VyNbNhdRWJPJoZ+iCfXl6Zli0heEKL1tK34aINsPYczje9zdAy8yCZpKivy+f+TJtTsEckFhnmrdK9f5LrEZSd255y75rVKQL2MKjrJSZKlM14i
UIQYrpTSVZxiz3J5rH2sM9o+DeYSqUna0ZnmpZMivTon0FN5IEY9eIcCJrtgPLzuc0t1q7Ew2gvYHm9WKAEPQugvC3R2GLp1uSzj7iV6A3TvE2x9KdrA+nTjXyN2og9Y
321FywZNVBspOC8EBzKvFJpeODyYWo0rB5BF5y367OXDAVEi4t0nOrEe04ujexFnIz5UyXPmhOz0s67qs7RcZoqrn1UukzlIQjaYziW4J047yyzaPMzK7J8VT0jUDmR+
SFvrOJkeHsrE3695mC82Bu3W5iufZM6wN+8aIXbsxUpOpN/iInaPoj/lEtrFKZx+n/klliVLMhZ5RiAytKoqtKdlMLFVHi9c7QVaGDoxGH4Af2J9k0nUFrHqqCRrLc1G
ylCphZhOMpFd0KUs0Hp349o+DeYSqUna0ZnmpZMivTpA1lR2Ndi92jov7EtFdjBYEe0PAOHPjMOVV4CI9U/PDu1cwduHnCc5zlJowt2wVNrCo/DkIkthRZZEqSbNeG7v
25jYwINSGHwaQhq2yohUJK7gooJLq7uqgapQwcwaAqSaXjg8mFqNKweQRect+uzlRoMWHoWKIyjbQl8YP81iE2O5O2UQZ2fLGU3hCLiAICZgve8ymNkD947ZoOaO/rwF
zNjkhvBBHRNcSm9Lm8PAyAB/Yn2TSdQWseqoJGstzUY88DblNTKZwwGmZnV4S0+aKWZToWAUKzEoU7qq7z0T52RJJY4rk7InR/dwo4V7KRAVxodKdfkrEFafbRt3Kyqn
FSz8qAwM4WCWd488R5/XklE6ad0baP3ZoUQWWdHqu7nwfJTni+sKBo/nXb1HAFQY/ef8LckCM5LbZZLZX6BZ9eOMzWBiEWyYB3Xr23WNM95qF0vczRG5kjYsQ30hxkde
lhss5iuY5HKXmyCHkLDOcAK2rtnQ+PjdZuVwryYiUTiZ+3iYK6EVQvsPqJNotL999WnwtzfZBhe0RJkNcbMUFFUiSHheRHfaUEecBpmAfRtglL4kK61UDzwfLwL1w559
sw5uAZS8W8XvesSy3wj7S9LUSQbCUfZXOQPOKfOn596Apjcc4q02He313LOLF1SEqb69r0DPBJKVsl0tyyrr9hq+EfAZ7a6D25O5Iqgs7DZVfemtbfLLBn1mXser+T7m
10+KIXsFYTOG6b0aut2atwUxxYtpR0JpBcxG+3yMtMTH7cWWtjqjHC2Y0vTybTd7VX3prW3yywZ9Zl7Hq/k+5mEW8yNkAhhGNQ/qptpaKgnJi9P2M7v05ohPcnPcEUb+
qpmqWKdJ9xKIn4qYuvwJbGUOnNp4kgSKP4AdyjX+YstysVFL4yHD8/9y53o9Y/Kh6ECzt0qK5fh55GIl9ERL/X8I9+xISbogcPwPZTEdNYo0GfWaP2Lww+jpEk8yo+sm
mD8KQ+aXmLk7OnpJrn1OJfHPVYrP61jKw5iBQGZbz4Xe+FoARkXxBqftGL78eBsuhH6pKV34ghuqqcnKtTq24vMyxxFeyPPbcmYxSkBUkhTr6yJ5z8/iKWumzgiz5XaY
5Bf6YO6RqheEYI8xx7OCrT4qns1pd0IOswGEt0rvs3GjAEFJs66v1YE0iW6ZjDj5dS7rhI4kT5ucgDA92PRYpvxe3ys/Z7A0Akzc0zSOQD/02n0BS1Jh7S0nSamh15e4
owBBSbOur9WBNIlumYw4+Z82z8mc4xvo/ifIQ1SuxU5t7grx43jnU1T+b+AKf9UVjtKvCIlQomGtJPQ7U69T17yiGRxXrXlgYBIwAIDIxd886FqwggdQG4R4i+tek5ve
dDjeyX2hgAkq8LGS2ZFHsd4Is3iKJJ/Bu5eUvG9titDu4TllfgH8y4Uxvw97rMCMnmFo83c8IazQxWNbcd6dvO1kZn8UwSFaPkMSTtF3IQQQiSzkvh5Gw/r3o4FAFGHB
I6hXTUvv6KBrCduTj7NNhvxgBlVLkI9DND+il2FFoZlkjb7owkbC60XvVJHOWzyUfcm2hG+IOPXPFN/6VeGMmYM803Tj+7QIo66Rb7AGcmWVfffLhyPV/314E4xbprSS
M5Qr3qtLzEHjxmPJFnLZ/6ROmJnmSMsXMDBbPW2w4O8rcsCD/y19AILYruzuCLQnGaB0vpPur5HIxDZzmLGp6wrwCIojb2bMKlbuMAO6+LBYBfRpKryN0+d9ih+Ddagd
gH8PhXYN/JALHOGN6bWoirYMzw/JelQOwKYe0PdIp+MemCu2QRj0cjM7dhYWeLMLXO7hHnk/duC2aVOtdfWehuT/ohkl0SN5+FwdXSNiFiBYBfRpKryN0+d9ih+Ddagd
I6hXTUvv6KBrCduTj7NNhjTJUpZhuWfiymzrldMFIuNvZz8WHCAWbvpxrKsuEkA/pHLuryMXFE/PRMjP2IrYZ9BzUDW6wAzFbGRMhw+I8wY57qRqmhxNdfnLS+SNexBy
2Z4h3MDRCDEjtBXMW2w3cKROmJnmSMsXMDBbPW2w4O99waJRCfwZ1vGTMGuwUfvtdE8GKi/68U0oc3PBrXaypEYzyqu69UgLQxJo4dvl9K/e9z1qrEwZ4WloQ1nK4n2A
LBqJ4f1pc07wM0ZTEOiarhi5rLu98kjo7dridm54hNvZFJEYVKbtccWGJl2WYCTts5+OhuOVHMsbR2HTDiKr2PkhF52BYwckfQ5GyWbYOr1rjkBAT4K9Fu0Qt/XM+emi
zJfCUQ1LLP6CCtygeBn1q0vBIBLse9AOzVQbP0+Ib8zSC77SyJmCm6nUDYygl8FladYOiL44xeboxF3TrS3dcaROmJnmSMsXMDBbPW2w4O99waJRCfwZ1vGTMGuwUfvt
z6fkDiEQAJskqilqMQzRCWLZEhaR1plDzfRfKPADeyrZ6fo9rCU55BGXqN+boeUQNl1E2cuGzVOtRfFC/qy4gWTJpIwpxkycGRJsy7JdEuaBrUD0CdsC0U3I7suLpnJE
Oz4VyjAcg9Zlj+cwFwFDXsYD/TYQ3k1/2JnXzvgEwb8n7fJ486C2XyZI1RANxlKKHQ87wozU++4tjaY5ADzpvEyLdslYY/o38K2pdFzrQ0OPku3lBRd92YBUx9asJzV0
iydldj7wohBhDviqq1KbUG4K85gWbeWyv2uewPJSEQqb2BNh55TQk+b8gwIF7NFpGJCKhVWPqWAsY4KpVwW9qGYs1XNv7ANxadjjWhu08mn5kziYotNPnbcFj30BaAyP
2suyFT0OyDthqmJaAr2uKY3oGX2WoIcl3ICyzmqh1r7TCRKwFpKlJTa7jdurrmk8BtzQii1v7F+UY+Anh/QKYRkFOmKOUfRrmUe255nnVsY+THZt4VvRujUmkCJqLQ+t
nkkB/8XjzUC8PGA7wwOAbXrivEeCHuXnLzQczth/yQGoHbAjKvjqZMIL7gex+Y5KXi9DwCX5Efn4BKmi2X9BjhspmTwWkSlG+mQNhmSGi6xi+rKOS4nrT1ESDN4p+Uzt
BtzQii1v7F+UY+Anh/QKYeznRYayb6F3/QQJA2NsewiWIKcKeAEbffmkAiA59CbmBtzQii1v7F+UY+Anh/QKYVDu7RlRnqU3+Yxw2iy+2rmJg53zh+uNLCqkG9aNimcM
rvcrB+LJ9cEo0RykI0HFH6wKQbvF3ILH/ORTcwzOjLyXfeV1ATqI3mxaMgZQJaUcCHI786yrDnnTnPYQoT+dznFTQ0gcvXqvk1d7T2wkure0U5GbQuPLHE98uUjgU8ot
we0YZ6urZ6dBhSChuHZ0Zgbc0Iotb+xflGPgJ4f0CmGKq59VLpM5SEI2mM4luCdO7aThxCSnf/ZWQ5129GqMTmTjwZHrTCzECRZLp2toLUGIWlWFAB8sE05iGr2aQwO+
ZMmkjCnGTJwZEmzLsl0S5sxY0Z6xKQoMmQUKIBaRXEL31lT0h3gqRiP6OdFLVZypIxMOkbNaNled8CcUn/JYQEcuQWL8VUWKOqV9t0cIJdd+Ag0NURNi8ehVA+0LePXh
MdtZRsQpSED7T6a2AC52MZNI5J/U61YElNV9enzXmJeu9ysH4sn1wSjRHKQjQcUfQNZUdjXYvdo6L+xLRXYwWI3oGX2WoIcl3ICyzmqh1r5BMMfjmAwiUjDwn6W0opPf
teupiZhgMeCVz2JNjwtYll5NYtPftNp4Eshx1Z9IC0MuiTSNXaqNLP2ngQTT08YcYM19dYvShFdh13e+CmA7OQP46AdDPFlw8sCY75GObAJrjkBAT4K9Fu0Qt/XM+emi
gJLt3efuJuTTUWMIhxVz+mSNvujCRsLrRe9Ukc5bPJQiQ/OI1nh49AH9U+sq5ZtkdJuBBBvZlSde3VhOTgDmf1kss7oO+/EvP3xsV6upIY4nskIoi4GGN/G/cCra0ovY
t4tonZ/uPsgF1gg/bcH8q6AJfqDUwp7ax+bSwk9NPz7KiCbRJr2HgYyrX3ljAm2ImIceTrhLxrBY62hwvBe2HYEvqKcS4kl6ZdpAiU0KllYYx9ey7ASKabKcQzhLn2GO
VfTzGeE6sjM6aEEWhcTrgwFeBog9tG9Hg70d094l4/8PgyAS1iPIJoBRVWtFSjIACGmWF+m/S3YCFnaEOhIradF9Rfk0m6jH0e8QTgjFU5Y8sLsF2kXrvRMRLxPusaYx
k7NgqW7A2QjmzqCt++YYCUpMpmug4DeThtMyVV/TEsRaisVmJnaffFJA45pNDUgQ+fKcRGxwySm8J9bh8on7O1rVlm5GSKMWuXx2WMuDXthgzX11i9KEV2HXd74KYDs5
A/joB0M8WXDywJjvkY5sAmuOQEBPgr0W7RC39cz56aKAku3d5+4m5NNRYwiHFXP6ZI2+6MJGwutF71SRzls8lCJD84jWeHj0Af1T6yrlm2R0m4EEG9mVJ17dWE5OAOZ/
Td+JyAOwzcqIutOdll3DguFuNyP4XcFCIBkp42pNAz8Q63ZJdBPsibXI91uvzeQEJaf62MZlAM7OHQCeKijr07Q2ltgqvl+i+/B2rqidkXUMrdAseR1zMhKpQmYQcUu6
UFNZe2lGDwebYmkcs8OZOu+r5Sj7RoMwg7w9fxb7adknMsUC/1sJidEX6BboozgSkLRn8p+TjhQAv7VQPDQlivsSxJjuG7olHOK5SW6VL6iAf02xD78ngwsxcPMmISa/
DY2F/f8NP1K+l4YO0BSVRlmphm9D7MFY4GNPO8pKLPqjhfrX02g9Ki8laRlRIxQzUq8lubAOLKSixGJjtBIL2QCK830aWWmMzNV0ysvlTNVStwSYKVk/24b6qxVbFnab
sbCxjhTGUxZPG4usDxQ8CGea9EK3fM9dZJuB4Wj65dQmm5Oi+XAhKKexM+yz/b3tAmpAurIMuXt/NvcTHzEXRH1T0OyRAe7HForXS7+5Tx0EUk8ynqSzJRbtgh8ZJFDr
n7OC/5/lqXTXS8RMx2JusBUE3ZTuGNhZgg15Fa2H4KpNvkI26lNx9yK0xguKqS/XREj49+JIHtYteSK7kvI2c8HnWE4PreWfNzPnHtfYwK5jckT6W6QNXwlFkF97sPSd
Oz4VyjAcg9Zlj+cwFwFDXph+0scvMkcdsIG2R/c2GN5Ppn9l5Aw4aC52FIsRpNYKRQwcurL1cOtuMPIRplEOEFXc2NxIsMKWfUqKXfZEP6QpQGl1wD9k+moe4aFzXIc1
NTi4IxQ3Cr2mSD4LDAbWfdrLshU9Dsg7YapiWgK9rimrCfD8QmzTy5e7SAhOnSo+CEh1UT/WP9ZIgziP3SlsnsYEKbvhLfKkFVq0vFBLAhRPpn9l5Aw4aC52FIsRpNYK
rH7lCAUSkUf2vonCiXtNXErBwAzcIsNAW2edsS3QbZ7tNo1TkrkT6bM6aISFW/4o43rfeZ25sU2LcTVwDmCeGWSNvujCRsLrRe9Ukc5bPJQiQ/OI1nh49AH9U+sq5Ztk
dJuBBBvZlSde3VhOTgDmf+QD1v/MjEPXlxb2KM2EzAI+I0zWPlMHWSZMRWYRZ204HmcEzAtP6wSVwuUCrOrzcATXVAjlkaqkVydCznPCophZ7iuc8+DBLkfBZTjL9nIL
VuOw95SQO/1Q7fKPYfQLnB297J3u0rmcogtdeZMhKqEUg5N7fiXKoPiWu0+/EV9LUXZ6XQYQetd9whoRPw9KSmo6EHrgSMwAdIoawpFPK9BHbE8R0jHvFGkRAPbPyPGB
85WpCuxNi8ySG2RcatrsxTlbDeb+qT9ezkFlH+0iTRAJ9qTHE3v59VxTgDc2Bxxpdq4JreCcD9yGADlG3GbPAubN41p7tYnYTfFm/pBc4zbRnLrcaW9UeZ9aPMIw27Xw
yogm0Sa9h4GMq195YwJtiJJoJCySArgci70452ehY9W6zNa+ajTIQDmiHSw7ic3fx83A+sMqbvd3e3jwmwIZyoQoEjBcGpdYgRznp76wyE1LAxajczm+X/6acRJMJ7v8
446U0qSuwAXeOpq8mDF/rxMObHPripb+WknCgZlG3F7ZH9GcCc9eAf/dJEEntS8Xgz1EabiWYqjL4YKML6lamaWEznYVm0kCg2RgavI5ICq1SJkjHqmwTCiiHFxtcfDj
MMrGeSMRvj/sNZBnRpre4aT/2CbiVJsFNzuUC6cmnaeLtykXsPHfZV3KEfSIGv2fwC/pr6VeUTyL6lb1jcHXBkfNoi6XmkJlHw3mTYTl4ZaI6fLzKKlLQqhOe3Q3rxOi
kExR3gUSWHkVpQMgV+0qJtbCSn7X5nEawRTkFFZpJ/vNk33nlxzUNeVxf8uD7ElDWEnNq16aRrR7oE41K8YYNYDS6Flqz37cVHcvMetLi2YdFLhb0Zle/b/etLohd4MQ
kSvDoLFvCHV1SWfK7bIzwYCRLCER7mBh4k+MHnlO64ljBjexLwjfnH8tdBbiJbNl6HjXIkucajMw1WzZoe91LmJu4OJ43r/pgsYnaHd3zJKE0PKcJM+wiD+pKAECTSUg
T/zMIU8keBf9Qd33EFDhkwrd2FFCMRhC1MXGkO3kPrqzdr+HDksYBIidRlQKjNeyeuYsyRojEq/8DF2CyR/+SSuU4r4zbiaW8IujtKjgvHxfF4bLajNh1FQYs7YvuYwf
HMqqxeItMf4DsmIL3gQFCHkA76+VFCYrkzMuXNkXKJSz6s4HvoNtgafnSWkCbwbAQDiPLdTn+um6cZCZs/M9GY6ZUy3qJDvXOQg+u2YC34bbwhGO/i/hrRukFVTM0i9+
ZBSflsvZkUsjtAgXFxEW9AHE7xfIMKKDCpigK7+ZtPBtIexqvVKue3w34uMG8ZGRnRu+6k9KS/9uQT10PQ6gcnyx2tTnFV7s2W32U4+lL7PCYfgj3ph+E062eWOFDemv
+fVdvE4ZDuFOMyA6znEX/ySblz/1p6HPZBlrKhNqObyBmt5pisEaLM1AgfyqQi6irmiKb28z6nh/zs/ApWR5V/y4PX4bja/GPovkcdJMR1GaVmOvBGNzOJFQ8VBCsQAU
1Kk7XRyXcGQKDmh/1I7vW3ttWlOLh/mL+n6y1O6geLBE1pcXe+6/avnnnqjrzBQfNvyK4lRdgFV5R1kYyNE1sZcf2OJLH7psfpZQXqA3M0bZE3xSU8yz1nU44YTAczpN
Jk9brZvsvZWxHH1CstKj6JR+zwmV8RArOgI1diZW9az8uD1+G42vxj6L5HHSTEdRnL6MrxCRAuFIUkAQ2hDipjfYO3Dvj81KtS0igMzAmzt7bVpTi4f5i/p+stTuoHiw
HZzLEina41/tOFyOQGriXuF/qRmqmMVLnWXgTqdnmCFOjNP/m4HNY5ALbNiXMpEoBMYe4ytNr92OL087syYw6ITviBlhFZU3wCBYzRICFZwBa3TCNYmuZchMvsNXmkk6
AsX5xNAIj8hqSJ9/7e0H2I8QT71txe53CDsAdux9N3ALJKH2DTh+2yyiQWjGtzgbdhnZ3HIuCccT9ZTxmeD5TeIDUiQxQtLxBafHvrr+FR97FyQFzf9yZJOT5VgF7ekF
pU9jG2s+QQG6k0tM+Gi0pyYOnjNYw/Ba1cxpwsOi1xDErrAkQcFvTfcc7pOTb/tzK2LfuTE3JJ+1AY/TY2c0pgByYGJ3rUWxSKRWkqkTXBqNcwT5ExRmJ0o2CM9dMmtQ
jMGRJzlB5bTr3zm7lFOiqkgsuK1nKYtzqMcrGPq2pCBM1CGr004SUAUvGghL0vCod48S1j8Xn+ILpF9PZ+1IqX7X18mzn9bQ/BvxOmXx32UJ3tLF4MewP7ACtC5qnKOt
OjhvQZ/VSVXb+8QttYbXQvsp2UUnhtKN1ID9wLqOsrqiPqLUJ1CRDvCaClvHzQni/ArxS/Z166l2bwIqCG9P+2KrTJrjigGZf8ZOg6zpjRnxnPW6qDnu20f2H5Lme9Ku
8b0qqSjGDgcV77iDxmUsdB5zexLkfUN4g8DnrrSflo9zvtNdWKRitceobBXNnTFYOkkOTpCZIsMxsHaNzbu71v8MolY+0V9FwcR+m/gQIU38CvFL9nXrqXZvAioIb0/7
BSnxw6CQ1uvcNmo4JIZTr0aTvENTnJz7Enu1pOtYzab2Dl43NsNYFOrWQkGsrVdKGSmnZaEplgwQoWy8u0rJLw622Tc3trDabLoqBC6qiXjGOEMAgTQVBzfSmz6WN/7G
zr0PpUFrGHIEKln0/UyEG7814/8ujryGmxjppS6vcddc87IOTcgLSaToZt+lYHjUb25K7s2f+U8YaM90W7c1wPsAO8567jJXE/UOo2mFgbiOMFDvk8QYIBnLjEBA8+5n
FOE4RApn0hcntkAaARytsRThOEQKZ9IXJ7ZAGgEcrbHVi9Hf4HRg8WL15JsjSGW5f1XmWeKMuMWfg7yuQhFDZKTrbhz59y0kcQCYD6i/6gNCpWC9afPHi/opedS5qp5T
5MVpeq2a2P8AiYZuiVxBqtlYAOiY4Xz9okTC9Kxv6KpILLitZymLc6jHKxj6tqQgsEqGr5FwNzh2VRv7OHmwmwZ5Bt8heDtR0yXvjobLKvoKngf0e2UwM1FJxrZu7ZCT
H/hOuJeSpRSqbQhZUTXAHDnaUgJhpmi7JLbIpK3FNR/pZ1xgPSj5z0NsMgV5RCwb2123uYmHK2mc8Y6AgcAsnCRXYDIGkxvmWshr5qfUkFcdDzvCjNT77i2NpjkAPOm8
H9IJ+I/WHrXBuI0a5/TgkGSNvujCRsLrRe9Ukc5bPJR1nWVsSfxAEKHStu/udlJXT6Z/ZeQMOGgudhSLEaTWCsnbDat/wj1oUstW8aODLOFZz1KO1+9Dg6+P9Wb1OJkt
3Ss0ARK8WLXZwJU/NeTu24BHWlRtqMZ0P315X0qBgIIuYpGIjaUi7tf3s84xauPr2Bfr1zHVVB2O3842R+Zy9gnsnXuqkDGMMgnEt5iDq7u0NpbYKr5fovvwdq6onZF1
LH9E85u5qmXdW4oMNxNsqrp6cIe3aCt0RWvxiwB0ndjtT5N13Q3l1I0DPur2uT4oTZ2h6QQyIgTjhf6B7tM4ycPUaeW6sxAeTsBWkX5AfX0yhlaQEubuEsz2BHCFsQfD
ouzq4bblBSop5j2pwpmvgFhQLQCHpR7x7PZy/qp4qQpXRxkAJ/LMvqKYrj8eA9XwTBJtBe/DsMcl5g0USSNtYGBeJDFK6t0ksyb5UF2l6fh/+88slzXlShTmGWrPrbFI
kYIoCuk8dV/+/54Ud4e8qA+46I0G7l0vzAiNjGNq8/W+9vpJt1i9tqHytlIvocKEiP7jVuaX46FY/B2KzP7BmkPxyR/IS9kQgzI32OL5Pio2NETnit9sy2UJFl1q+zV9
OWhWRavz53D0a7HZ+7oa2OzGta3236BxrcSeG1ky3JAX6Ml7+BZS4N7c41qTW+jSFRe1djX0pHM7Z4j4Xv6FvpsElhNgON15aDVlG6I4GCQsf1RKNVg0pBWlVWn21EtU
+J9h+KovGBMCYQa/Mj5O9/4SrKyeYFTCWiS0VAXXfmDLvdoAYyPZ+IO/lk+TW2T+a45AQE+CvRbtELf1zPnpopmpe1gDXeE5jz3jUudqJD1V3NjcSLDCln1Kil32RD+k
zc6q9uiwWQAz+ylDVCtFslpb6VbQr5LuLiUFH01P5U57k2x/lZfmsSlOaWtBaMX5qFyo268r6To2SLoSlT8WmlNjJN6tcHSy7WNhxKUn2CLfql9fgt3f8oNFGv7sTvy5
4Sfxrac6YRBBS8u/9JwWfay7AieKG2XhjDpp8/u2lNe5BTTcNMRKvuI63vzxvYqPGpVkP/0O2gcbddPaIlTj00AQ5jbiwiRixlMvzCK8kkTiKh2rKumQrmCEsOw0jezu
Esx/MB2KVACyk0R+ifxZVIm5jBrA+x2DgfUKOQTcuKb9IOSKqQ07Ww/E2zD16Vr+m9gTYeeU0JPm/IMCBezRaTmT6dttjlylPof8UIFiUHlfKzomxJ1htltGnRRtNUv4
r0mQHdh0R2xKLQw5P1z2Dvy90IJN4gVJkfg0kxu1G5T31lT0h3gqRiP6OdFLVZypt50h3YbP+u9syWuxY4+VmpUl2fJT8Ot7wRMN2b+G/5vVzcWQwwlSiWPJw5vnsxIr
SiBrMzsvSgjnjzp5z6xQ0YsnZXY+8KIQYQ74qqtSm1B97v6ztoQHZYjofUKcxSJwT6Z/ZeQMOGgudhSLEaTWClPPSxBcfcxVu1XdxnPQeUo+/5fsfmzELLNKRpit8mR2
MVV44SUIULWE19DUWq7XKZCf7b/l97s8kwm9VvlSvJGuo56jhlYN4Df0w5V9jkIny97AUiHM/DkdT02yVCIvloC4l5/CQ2h8nArGpQhZxZXI5lam4UvfsoAoOMUpGUiU
EIks5L4eRsP696OBQBRhwSDD4zDS+UHhCedWPlxVBGb8BjoScWxpbiQf4sVjTP+LiOaAGLHBYLQOWRd0k/mDFh0PO8KM1PvuLY2mOQA86bzct+EImtcuJVLMUD5XPuHA
qVu6MnaBCMysuW8+bF32tJCXtHUbvcnUrHQDnnoZso4KZk5IfTF5am+uacEeLSodov7ywEBicN5gAXl0VWOyEkwwb5L46pKBAHhEjheqAkbjT/Ns5DLd2P1YArd+ZEun
k2h19JglIHlEQD7KreUyrt7SB6SME9CU/ZXpv8AkDTRQ4UnBkDIrATBm7se0jqV8IsvDEyu1b2gMeluIeSJ/ZmNo4F9EfKo24ytK70pUIdjLTQKawyhWTq0qzQZ12mUb
w/W6SBrSGGb4M4TJ2SnbwhWp8Logo3lVQP2nJWLnQ+HHv/hvY0Ii5kQp46pw3Pejdwoc55r/ehbabGiNxwMhlE+mf2XkDDhoLnYUixGk1goYACG4zY2L2h/IN9NrIY8u
tz2cm6BQPJD8a2YttOFjBzkJ/s9u7Gk7H+f7wRicrMb1mfcSMNz0h2XMpzX2Xs//LSmtpts3zMF1qApAF06rPc3OqvbosFkAM/spQ1QrRbJdsCZx6vK/96gPqsDxak7C
mva9vr4JiUwo0pf8Ttz3uSDa47MapGZVK3gKUfSgItMrdD0UjviTO8umh0gr96YlBKtM4dLVHmZlqLRtQomxkWYxqMN4BAsmV9BV9elA71FvZz8WHCAWbvpxrKsuEkA/
lw+ObQ8GsyrQhCMGfkmrBqan16kqYY0FGaUmYx+MoH2LJ2V2PvCiEGEO+KqrUptQ6ceMPsBYUdICm4eOvwvsxmTnw29GDmZcozuLu5lWZzbyav7Lk6e3IFACMt14mh4u
Na0rRCPKuzNleW7wB1iup5k4w6fknIt63IREKmAVaoH7j0PBEMk2P8v9GizxMvkFuFcItAMubko5A3PjdiUz6Z5haPN3PCGs0MVjW3HenbwKdPjK8+hCuoC1YCZ8sNqW
T6Z/ZeQMOGgudhSLEaTWChgAIbjNjYvaH8g302shjy5cQ0P/+qQc9Zll0CUSnhLyGr69BUVQlXIVeJaZZKOqvqlJ+2aYK2JEbxcc2ku3y4Gb2BNh55TQk+b8gwIF7NFp
8ocIslvyfjCKfzz2D2biXjO+gwYKZqlMGE+pzH5Iy2kdDzvCjNT77i2NpjkAPOm8m7bzTQF5LNaeX/g23Si23ZvYE2HnlNCT5vyDAgXs0WkxwNytL+sYSrTWCKnZibFW
vWRUKqVhFhkLTv/mXkgUTitFA9X1IU248F86qtWRXeYpq7c9DrjNbfsn1mofbMFQyogm0Sa9h4GMq195YwJtiG8TOkxHHaarvkVsyxNbJMsDoS9BbNldGAoAWmlDs9BO
OWt/aFcJU3XMQlu7Yg11TOy75dGAZ1iu6WPuZtfT5j/e2DfolkiNM3wPtVD1H9Wyi/OxW6RoZro3XIf5QSmptR5nBMwLT+sElcLlAqzq83BlW01aUONYhMCgq2Y6pcJ8
PzzzzxFlQMBWFeiF7OS0r5jMhgTUF2P6jojFwL5rDN0PJMVkT6SgGrUlUbEYwLM/PzzzzxFlQMBWFeiF7OS0r1tBwR1u0P1OujIqJ7g+lirj/bkc1BJx03iblosxIkFM
of2SEnUt371Ks7aMnHIzprX0KNpuupEyuj1x00UmrMjz1zWvsVGhDEyekfrvLQ/jT4o+ycFjNLai+e5fFZWDzwnr3aCTBSePlvSssvOESjvsAF300tmjyI+L2k444QJ2
gKY3HOKtNh3t9dyzixdUhITeC0hgYM2ANwGqrx42AyPE9jvV190VI6vQ9us4gBWxi2hPnUSP4MQ8v60wkXjCJt87eGsX6gYkvacBj9HvdZE+EVjclhk5GMVNqGoHM7qC
8nNOH25m2cie5+yIWMRR7tYktEUR6+2QJWBl2C/uZcuGAJRjUWJ/zlrYexbxJxF2aBRKWnTzIEaGy9yO+1VgWjxRlzPtDEE73Zjg+cOFO0AJPtnJgZfXknDdNjvd3cwQ
IpE+Zun7hl6cJcc9JO7e1T8ZNTojtb8Do2OcPeNKZwePZrCjTIO+Q+vW6P+V9mJq6fit4C6377VOu20aDweELz/aqxE+nhezx+L6LFdldSfYGm1OjqdqN1T4JJrmdQPb
a1WcsKHYaDTx+M+18fuabk8Woa3vCUibEu9EBQGxg62ii6bAVrvDv2smY3SbaEo1YL3vMpjZA/eO2aDmjv68BXYVFXW8Ph0+MM7ygckdEfKiBz8lzWwRF0ggCzkL9Q75
vxlnUZQTQdaZH3sh4+EurO3JSw4kPcJLzlrtLMiwITuCBi0l7v+3QlUvf36tFf7Uv+7+n1uFONHDClOM3nrtdobzF25e54946bpCf4TzGugNPYo6uxP2CPH3Cj26adE/
Txahre8JSJsS70QFAbGDraKHpbFxny5DovaT2BmrkSxTYyTerXB0su1jYcSlJ9giTJO2jrOfAJAEu8OA+wNJc+HOobfzxpookYwTe2bwPreJgjVFapPhtt2F3ptJ+jtW
nKJupSRUkomO2eN0NVgPHZFca0DiazmbKzbX2pIzjhnHFIB5SnOQNwEg+GhN1gK/S1I694rqF1Cy9QeUWA9dXQo6ntuzwnL1ITawu3lwToa7TrzDufa1QwAZOHUzK2R2
41FnfCeZkFJmaJwalVa5hKt5CyrlZusFMLPsXxFiXOSL9Cc7PyDE4nqTgZjDyP6QGUyhTz7s7mCobUZGZNbpgmCUd21aS+PKR+qTxdQmFi4J692gkwUnj5b0rLLzhEo7
DYNsnSXTYY5S3BjV1BTk5XLD61xHv+ffRNZQxfXwHjPdM30hb5jEKszeFKSi7H9ZjuR+xMHz0DBKjvSMagaI/EbQClGMsJ3g+BoXMRtM1e4SOiJRNUvH0C8AcO4G2tXA
Na5CYMdrJ7f1BfzDWBRAGDdeI56snSwAESCitUKmTl3ULq04smv+ZwqDydshQXmtNBlX0T0Fb12NVKzc3NXgijdeI56snSwAESCitUKmTl3LZmY4F4tvZ2ljmQZkbOPu
vY+G/tlsq0KW06KZrjICurUb85QR0xpE9zM44JG8SD7AiBnAsmPMvEVlX2Tt/WCvWNxtuqErKPhxJdXOZqDkMCc9TI8VVfxwqk77JJv5rcjKDPCXgOaxzteBILbK9AaT
X6M7YLmOsKBbLwy9DEq8QsqIJtEmvYeBjKtfeWMCbYgysuJBeuYXjsG8Pxu/RCrqLyAFnLQrQDhbvS3+nJra0jFiZ/1N++J5mriLX7iVoF6u+rvb7jZvRQCfSzvVedF0
yogm0Sa9h4GMq195YwJtiAM5rBUtNWy9qnDszVKYb35+6dmKoT3Ebkvvx1SQChwhyogm0Sa9h4GMq195YwJtiAM5rBUtNWy9qnDszVKYb37pYScsEhesrPAFeTuogfbW
lkfiVouvsklfgOyR/fbyHgM5rBUtNWy9qnDszVKYb36yYIjxReeoxGGZ84CgYjgpYpFSLKxqZHuHilqlccSaMWR7iWcHRe7i5c2KGOJTZYqynE9KyWHQ+VlxlSAuMpTU
igZSiMPpHqQPq7NQSccZ3euIgHYmJts0u6ITD2Einzi9JP5xZLRntcDfKWPcx9OzrsgnB9zSjYueDo1mIF04OXSFhujwopI6nXIuq9R+qXpDQCQb9MAG4UE9hkQjIOIP
kH+R5iaAROlsVfKBgS07aldX7saD5tT6bsPnQCdox3cmnXdp/gLNEPyYCh0GjKel4h49K08aGem0bm/AE6/r5tIl85pMPMM/ejdTIr7LJceQ3U9q3FAufoBEPwYYR/v1
xib6v2ng652CKMKOfcWkqN7YN+iWSI0zfA+1UPUf1bKqW601lxVVDNQ4/GTl4x4Fzc6q9uiwWQAz+ylDVCtFssm5/9e/gu0skg814E3EgDriHj0rTxoZ6bRub8ATr+vm
4zNqPiBp3rP1JYdLTbj732n3H9NWKR01H4XUpIQcRJgxhPf5IAbowPSgd1oDX7PvvbWNJY6eTH4cqDRKSZ2uQNKGyqdZT5TBl05zsFnDwLkQ5zZNCHEHVkm3EYAI/cl4
MWJn/U374nmauItfuJWgXhObxO7p54fZPMAi+t6A48CXMCDc25OiN1PjAaUxfcObPGnDdz7yZBhlZEZ79oomFTVCCxzgmNxwXxO/0aNEU2p7FjKR7FxAyyuafiXlw+UK
zwL9oEM5mybydtbqSNOBiE728kUeZ7sin9oWLIVFvlPbecdCX43zBQ5bcwDv6GAQCjAajx/YYi5jqQhDZS6lcAhxesbW3y39choPQkkfK5ZSrGHc9Dheh9P4P5GguUzY
0WKC3++oe1lxyYvdh0oDY+44V9XJAjB0WQqKvSBHInzsaF4lmr1nUbIDRtywY/gOHeRTWWeUq1UwPd5hrCcgf3dScausXeJ5hGascCe5vrQqkVG98WQv/ozHexdktIC8
p2qcmnoHiWdM8d1vaqCWU2C97zKY2QP3jtmg5o7+vAVXWY8aki9edQhsILRBN0GgB9msefxLXvUtIHVBlRVBMbIFNhX4fE0iGrgbx+h9IiWAh7kAnc1r3kTTiDdxk3hN
Fv0fLzIYznIXsh4WG3MdvsJ4aVU78MKCa/37RhMQ4hN1ixs9Y+Kx7k6oYsl5RhWm9ofghizXJk2//Nh4p/HjeVckkC5TdoSyINSPJsWb4y5/28iMwTVqnZ6rk6imyAg8
wwFRIuLdJzqxHtOLo3sRZ4vKvqUAxMn1Yx/4GLU9PJXcuuR/morlsLM21h610D6clzAg3NuTojdT4wGlMX3Dm6rMxB7T8oZSKJ3kwyGrex2DGEGvQeM3QGRgbMspUSII
7Hb+B2l0QNnTWMM2g4VRmGc4pa72nWUGQh7HH2zGPRj4olUzT5ombdI1SbsmTTeSXm/isratoKhldbZTBfLHnysv78eLjGPJjPHZxpsB2ygPJn96Fxr7rt7ZrLcbKE/R
oWTldAS3QCQi0zc+gm/kC4l3YNcqp1dfw6l5rgQXh66pGghEgvQmbaNga6KdHtgKe/1zOKUQVlQKiddrP8BSu3/byIzBNWqdnquTqKbICDzdnFF/pAXdg6FdAIyt1HS9
KkHTYLZ3eFVgR6Fcq8b8rHj3UYY0S0+Yk7uJahVbTBPj/bkc1BJx03iblosxIkFMN14jnqydLAARIKK1QqZOXbbng0xtNnld/dSELjm7j6mMrSyyOCepCIwbNfBJrywp
bhHaejfzOsXC5TexcSMQkkz0pmWrQw+H8R84rf67P4fexGbntnWevNmJkPVL/AUy3o1+5jey2sfGJ+5jpmlZvulnTRD0fTKKcMe9gW90IVPjIW+L6/aZ/r4KuyW5BY9U
oRD71yvPU7mvtU6oImrYYYk1BYlHMTZ3B3Fk9q/jvA5AskAKBWoPhjhy1doiv6TbQBDmNuLCJGLGUy/MIrySRLuT5Fu+BgACp+UA6C+bLtJZw+3zqqmSBR+zPZ1Kz6zx
CdHI99/cGPFE38MkQv7X5zytD8f4KHDoyaK1cn3UWwLxis1MERajAdxLqcFysLVnyogm0Sa9h4GMq195YwJtiPUH8hdi6dgDciheUbyvzbjKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKqxEYc4ZTIt+jh3I1MQDsrQsVKQRByGDQIIrBrQWW+c6skKh+D3K3YJSN8zpkS7pT4JPtnJgZfXknDdNjvd3cwQ
rET20/yPopKiffaDmGE1+cqIJtEmvYeBjKtfeWMCbYiJr1+Y0WAaMj/ktP30L3Ua+5oX41spF3D8p80leswsLSG8E+/izOgDZtCcT6SY28Rgq1WQ1al/4sEkvWSq9JaG
1/t95s0mrzrugeNvizufGcqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IVOnKOtP+caPjsSiR3xSqHXfv5bUTR8gyihYzKekp8rJgDITO7hq5vBc1sZU8qQIM
PDSEiXhe7tjEHe8tsX0xVv5Y0IrBpttDMmPH6IkfPmh6zUp2SlaE21s+qOovTy/4T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCDZBCVr9VfGh/KGPVTGrEM9
y8ShwbbL09ZY7UAE8b0WSqfuasrOZKKFfKCUbFAiB8GSgwHaf2C/XgXHxwdvTiMOlmJwqSxzcxgAuF0utn7RHvXgIbG2KXL7lT6fOiJjyKp9fYBAWXKLMO9Zn3/M03yX
3FwpB767aQ0GHP8+04s+2pZemkoHXWOktTry+ZmtV/AzlCveq0vMQePGY8kWctn/99asvlT8I0Rakyes9mh2McqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
+5oX41spF3D8p80leswsLeGyB4FFotbluXPSe/r51qhgq1WQ1al/4sEkvWSq9JaGrLsCJ4obZeGMOmnz+7aU17rPT6X6LpkLYO3q+7YpOVzKiCbRJr2HgYyrX3ljAm2I
VOnKOtP+caPjsSiR3xSqHXfv5bUTR8gyihYzKekp8rJued75yJMlPYATqw/hR2yWPDSEiXhe7tjEHe8tsX0xVrTZBNV28cHZekQcnu3TyquUt4nhQ4Mu4PY+rZfvVABF
T0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCDZBCVr9VfGh/KGPVTGrEM92bPoOpfcTwbFb0FbraCaiqfuasrOZKKFfKCUbFAiB8EZIHR6gEddMQcEoVU0LSlm
+wDWvearcAqIUiKTI5x9fvXgIbG2KXL7lT6fOiJjyKotOAzdk3Fu0STcvCDdr17U3fdyYNKT1Io2V6H63wgKockKh+D3K3YJSN8zpkS7pT4JPtnJgZfXknDdNjvd3cwQ
rsSlqw/tvB2afNIBAwsMfsqIJtEmvYeBjKtfeWMCbYiJr1+Y0WAaMj/ktP30L3UaBbNl57kaeVZ3SFrFpfQa1tiMYD8eF9P3gXRMPHskkYiXAHuuKShezYjls0vGFEp5
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IVOnKOtP+caPjsSiR3xSqHT/aqxE+nhezx+L6LFdldSdUnYDYG99HjGn10FyEDSBc
IRj638TjUSFFWvykHyG0UpcbJgrK8gqtte4y63U3BYFA/Jv18/j4EB6RI1o14dpXT0AdSo0+Ioxd3pOapgecMTwTKEgPkf+G3npp/y9Z6oWSJTVfIBkgo1pThGGEXjTG
VE8UNg3NkkHs5eb0lm1z9t3bk7eB0B79tYM6g1lcSjSii6bAVrvDv2smY3SbaEo1U2Mk3q1wdLLtY2HEpSfYIhWUlOWGomcVSpgfSAS//sAtOAzdk3Fu0STcvCDdr17U
Uom29Wf4IgT3tFDKK7hWXGBgC+xNIFxLAhtED8lTcGUJPtnJgZfXknDdNjvd3cwQIpE+Zun7hl6cJcc9JO7e1ZDF+xfu4ZNyscJBSqfM92A54assiAOsTvfX+GH4ef2E
ui3vuQ4ZjxyD8YTXuFEPEAowGo8f2GIuY6kIQ2UupXDNpDa50ckJAQMzdo5WTPDF1iS0RRHr7ZAlYGXYL+5ly4YAlGNRYn/OWth7FvEnEXYWzehi8upxbgAPaVhV8n/e
HnxxE58x7qzsr23/eeD5yj/aqxE+nhezx+L6LFdldScpjNm6XzNVCX2Vq1aO/ENuIRj638TjUSFFWvykHyG0UpcbJgrK8gqtte4y63U3BYErL+/Hi4xjyYzx2cabAdso
uuajdb7aPI3ezmuDwnVNSTwTKEgPkf+G3npp/y9Z6oWSJTVfIBkgo1pThGGEXjTG+TsQj9TWLita60XlReCw7N3bk7eB0B79tYM6g1lcSjSii6bAVrvDv2smY3SbaEo1
LP+fkGk1qObC/MHRAAOxW6EHcjD6T2qzDb+PN+6O61ktOAzdk3Fu0STcvCDdr17UUom29Wf4IgT3tFDKK7hWXKgdpdaTfu+hH93nCkY+iTgJPtnJgZfXknDdNjvd3cwQ
IpE+Zun7hl6cJcc9JO7e1RydVznxAXW4d65alpi5LOUVbFkgok+jdTwUlyJQItCV5Ni7ILyKbh6I4QB6WO8k/k1/dFQI+bNoTdA3CtXKYvT3YcnxLj+BZEuTPcc5ryqF
1iS0RRHr7ZAlYGXYL+5ly3lF3J890MeVE7UULObyetTKiCbRJr2HgYyrX3ljAm2IHnxxE58x7qzsr23/eeD5yuugJK3xwb1piENrZMCfy/LKiCbRJr2HgYyrX3ljAm2I
Figv/smMwiuSygu3ZXr2LcqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCDb6g1CQTsPhEUzii15lJt2
yogm0Sa9h4GMq195YwJtiN3bk7eB0B79tYM6g1lcSjSih6WxcZ8uQ6L2k9gZq5EsIbwT7+LM6ANm0JxPpJjbxDZlloNdhddpYOAaTVdVPMdnnprIR08r0t4RSPUEO/eX
Uom29Wf4IgT3tFDKK7hWXCYMo7bBXL49tfVn0pTcvjEJPtnJgZfXknDdNjvd3cwQIuB/07MIQyWMhqcb95ufYGAMhM7uGrm8FzWxlTypAgyJr1+Y0WAaMj/ktP30L3Ua
rEy5/Q7pvSjp3g0+TBQk8o/m+CTyK1uIXUUyFuccmJ6KmmltS0WtQRnAdf8Epji21iS0RRHr7ZAlYGXYL+5ly9EL2wdvNL/TOVyQyufUzA7lj+5Qxbdh+IpduD6hqTcq
HnxxE58x7qzsr23/eeD5ykTb0PckcayTEhQPYxa4EfATut12iiC0H2gb/wcsJLunIRj638TjUSFFWvykHyG0UomCNUVqk+G23YXem0n6O1bcXCkHvrtpDQYc/z7Tiz7a
r4Cl9BpgM63ymo13P50LVTwTKEgPkf+G3npp/y9Z6oW7mzkS3og1g1UH8BSLEXfEeUpGe/zsrGHBwlmYozEG3t3bk7eB0B79tYM6g1lcSjSih6WxcZ8uQ6L2k9gZq5Es
zh9hRwtv9+sm/txsWiWsqR8z9roRAmGHV4cMwX5vCKVnnprIR08r0t4RSPUEO/eXUom29Wf4IgT3tFDKK7hWXLhcGm7szcJaKl+yKzyRPJIJPtnJgZfXknDdNjvd3cwQ
IuB/07MIQyWMhqcb95ufYC3+LVS+fm2nX2eWQwyy0yj0ysJc478Ct9ErenMeavNJrEy5/Q7pvSjp3g0+TBQk8n/sDkRg/CvyAFo692+Q1ueogDRTURuwWo8EsG90Pt2s
1iS0RRHr7ZAlYGXYL+5ly9EL2wdvNL/TOVyQyufUzA5bQtbEx0pSk4+HSIGt1s3jOSD3RRTiMWmcUg32dpP+7EwAmsMeYpW4YWfGoZsD/WnKiCbRJr2HgYyrX3ljAm2I
ZrcLGKwLi1HmpNbySNKCssqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IT0AdSo0+Ioxd3pOapgecMWFNnfnyFcgmOOvBDq22UkQwzRQ/IEAu6lPvglUzIp4s
yogm0Sa9h4GMq195YwJtiI8ZXQLQemNcvk46DbU8sD/KiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiJQcVJWN3VgEeoqzEzbIFtG9045czkV2eCTNlsrGTLCI
BkwGUKIWXrK+dktXFEs0hF6sYDOyL3zbXWpKIzZRTGDamiMzxohJX9QtJGphnR0Uk2rvUTOd0G00kj4PxSgxpg9Rw/+S5UHfjJdWkfIeInSiRM7SttwMGsnPe9/OG7jd
yogm0Sa9h4GMq195YwJtiKBTe4B3k/mbHjIUfqo67SJAbdMM6xByhn5G508Uj1sF2IxgPx4X0/eBdEw8eySRiJoakQaIEjpQrWyiJppKoJaTqBrmQOCIctpiRO8Im3Jp
0yGRnPZE1s62DA8g752IHPRtryrgih5z6Xf87FCiV1aO2emTXJ3IUtJlFzayC1SL9Imwij6nEItz1KPL77uvMM3CXs9DpngQRQY5VLoHf7nKiCbRJr2HgYyrX3ljAm2I
d+FUBXZ3L3OKxqh0id+YDKGhBBibOkZYDkL5Wc3evRTrGCiEa1n5FRCgSaW8MEXKe21aQPqY6WRt6NIhxQH27Np8KaxIxCfwRJJPZaJ4Eil9SChKNknSZ8s69N+tqhXO
gnOzlbhy1j959VH45Izi9MqIJtEmvYeBjKtfeWMCbYgNHbaqvQlTYDBMSDdWQGuUyogm0Sa9h4GMq195YwJtiHIHLql8/FShcQ41SVHzY3YfireNt780alpywnxKv7es
V7XU5yxqC5VTGaaaZ9W0MGnFc5W8K+JgXR/hi7QeaIx3KxmAGr9BoVcuPk8HgRDBw3tEl73LMKk+Cn0/9r56zIUc5zAXPCFOpd5czvGFIhS04dGMyIsfMTY6+Nez3VU6
ZBW6B8WbMtfByuI0e1tCQGYbHLL0kuhae6i7pENgo//KiCbRJr2HgYyrX3ljAm2IKbAWmvuvd8ilV1icDV9dy5cal+XwjuLW/Ad21xRK7vjKiCbRJr2HgYyrX3ljAm2I
wOvgWrm0GzTcxJE0ZMdWwWHggyG3st4ZUSovnxIz1EWDcRdOfnzDCIY08vsxLu17m1tIG3EDi96Vx+TYHOsfoMqIJtEmvYeBjKtfeWMCbYiqZNYNfjRSzihQ8Nw8imlU
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYiqBo+TDdha2w0Bhh+sXXRLN3OcLkli9FN31vnndyclVuzHCAZyEzPxVLePXtMm18/J8PgCLzYC/VqdgpdS9Wsv
yogm0Sa9h4GMq195YwJtiPEnmZ010YJq+bt6S6JgYT5IN2Uz6Pxg2+hgtk5u141slaz6DvRgTEG2Ci4i7xdHEYNC8L+R3Rw2EovIl8X/gx24qrQZDcwWujDcuwR+FUoV
d1Aj/m9bekAQO0ntSgY8A6XtOaJMxrlulq4hY4/uHOZHFuovdJtP9FKfvqvAwGo9/iRO7HScw315f4DcAW5iLY4hEQ/vysWamWXabndot/bWaLJ3z3eTjJTLOZZ1xDRw
FWHJu2CDQZH3vAxztQoGjblJn++I2nr34CUDxN/37bvXfwmavFUpEoZQfYCyzAS6peMOb0s2Jf6fGzmn/LKBt20z4N9wXwPbXUURU7aWb4LeqvKtvW/cHbDaTSZHAHEG
5P+iGSXRI3n4XB1dI2IWIGDVTXo/DA4eN+3LiqoVNZ9hoF5v+hKm16dSfudZnMogt0GKUG3QeSD1BvqQcQntkNryCTTH7enMesNS1WCtttylUZwQ9tF9L69bzWMaD1fU
WUIPlffrjfFrZ0xZPMqonafsbYvX6AGXwWfk3BbwyNpM/7aMejMOa6VGMlf+gmMYKEKqQyZraYXuXWBx7u+IRRu033Iqp2OLCct8GF6oNZms362if07z3/e7E36v8pH9
yyxdbXe1k9M3Q3bFjsahKM1+qYxEMYqeC+WFmAW9sg5MRnvxqbFGdq+uMv2EpgpckYmG/rMM6dc1YHwwSoa8XBupYkQsCNYZCYMiURVevf7OzsaEbwuumwjaWZ4lJS1u
Ku3qQQtJi5Tjk/k3i0WpXsomlX6BkPS9k6d+daepqaAFxaPNGm0UGyyxvPP9Faz7qAiFsBwMgBtoaRm3YtERUxF15l1C8Cma1b0JOpinkUjWaLJ3z3eTjJTLOZZ1xDRw
5WcsWiMeGIi3Ic6Nt7YaOrDpxRc5Ot38BslOec+mw7loEeFlKFnCnj6gJ9lQ/dTLLVwsJd8/eKygab/o2w5qTyI4p35t/8dL7EuGIX925jK5Ddzq3FFGVjsmoN6eSw2O
qgNhB9I0Kh7O+qvxs+q2Rl/QkDXKlbhEoIit1MJivrr45tcFdEVoxa+PoVmTxCDqBcWjzRptFBsssbzz/RWs+8L7fDgwyi3tnQLsMcLpUXKTHuQ270SXyMPGzqi7UICm
XPOyDk3IC0mk6GbfpWB41Au3Xq2kKv6D7XlRulaz4k9h17CzDs92XadJHtD9YKMLCZAWdNaBlxEX8Onz1P7GIIq763yxtgAMa5rd7Me+ez3oXbU0QSK9GDeCBReutNPu
m8SLA5ONnzEw+jDJGbKvamD0sMBrnH95pQZXDrDkI/rQLHtHMhrq3yNQmfwKtjMJ0POyg+6mFaQ/GvHYETnt2iTUa49Q8m2nuM7PD5fPW2+i345vcQ2Z68oeF2BiPbkf
yxYGwLnnk39oMOJtjGCR2EAbhQa6IvlT+Hvti9Da5C2F81oS06f5hl9jLzgvj8TQegsxR/DX3rWN0agLpPLKLdwftTxlaP2xAtPr4TtIFgMzlCveq0vMQePGY8kWctn/
r9x07ZvInyqm9h/GjqXhX06N+BuE/ktboqe3KtYePZunam4zAepcv1j+g6WLj8wgIwmr7k7tisq0p2E//OKUxDihw2A97PaxTt61j++NuPAE507xgj5PdOf2/8xTrPzM
6b4vaFjMPSBDE3NIUNnXKUe4j+4TyuPkWrdVuzKvOo3uGUOcLQXO4oC9Qo5DzoGvuKppEgO64QpVx1Kbbbif6Sa7DpzFRl5WEYj4n7V9kctIAwVYRdGnUTGVuRQt73DH
6NF6Mf49FZqe0n6Xi+AmS6LAkqrN66K0QmEbaFAB2P87qbGACYWCEYVD9qeG3JAXK6Kh2pKDJiA4Rsm5wbL3xwmbzPExbhQpAgTRi/SqjyDMs5b7nKvQm4lf8gacjbv5
PAEZBMsPd0FnODZQLbduBByd/Cve9cGXPNrRmc8jKuigoMmGpNfeTIgfjNqWk8SHek2aCPSv+Fo6K0MZEG8rMVqtKJizja5DdU1RerzhPLKw27DseU4sD37CTI6D63v5
HL75EhoHB5eW5vXYt9vzDEuLKkToCnCRF5Wy3sjfDsEBlLMVHxunHg99DNlWxVsefmfeWVBuhI7ZiOgTQ1zitNiV9jIGbcfAQIi2C4M8FbdbYgHJC/40jl5QfhuN9OOj
21oJrCJe0/Si1tfGHy4fu2OrnO9WuOFv6fDwnwaaRieOiV6cnbR76W6EYCmObvu9lxsmCsryCq217jLrdTcFgTbea50g17+FvfnWBIc+iAvkRovbOwM0qNa8D4G8L+Uu
cRHTB951Vq+bq+CU6vR4zPaCMrBi8SaclIr3AfZ05j2LaE+dRI/gxDy/rTCReMImoRD71yvPU7mvtU6oImrYYazl8GfOGYBF4LhGst3ms7gd5FNZZ5SrVTA93mGsJyB/
IT2bmFacnZbQps4mng7+Q+n4reAut++1TrttGg8HhC8/2qsRPp4Xs8fi+ixXZXUnCvAIiiNvZswqVu4wA7r4sEscRUUp4vff+xEC97xgudfRYoLf76h7WXHJi92HSgNj
TuWytn3MpnEcC+cOQBA6DUtSOveK6hdQsvUHlFgPXV0CxC9XtFYWwAXUc/2obhMxemqE6+X94cEoXB6TJqEjIuRGi9s7AzSo1rwPgbwv5S6+nmweBpge5aeJStryyIsH
BQBqanZRk3LSMsx4FprzMoKWQUszSgTV3K2lhiUTnSfR7RMI+0jihq7aIhZD+06+SxxFRSni99/7EQL3vGC519Figt/vqHtZccmL3YdKA2N4ZRj3yeIw2hgigMqYZAJp
pwsKXroggy6i2++gxG1ewOch+xtdBRQtczVnFSAzdJO62ge4aXw5b937mKou5IBvY6uc71a44W/p8PCfBppGJ92cUX+kBd2DoV0AjK3UdL29QShRXX+M4NJ/kGL+USwy
ooumwFa7w79rJmN0m2hKNWC97zKY2QP3jtmg5o7+vAVWyCYaU4mJkJJ5tszcE+UkM+08jMsWX0fH9BKiTkzaIbpIuJfO1bormDO9/rwAlVVIAwVYRdGnUTGVuRQt73DH
BJhiWD4l0ker1E/8667aj5ax7QhRNMJRFak68J48Buzi3ycuWfrLN5IY/4MIyGeT8AxPHfjynPXC7Gh6EPS44dDEj869zF5rMBOp/Y5qptPzLJup3x/2Z+xjdyymrXEE
53E9STuMZYpgiqjknZPUiyfEvH0MaKuGgrVHzhHXWUYVPEvHrwdImTHOBtiQwKr7zszn0XJmLOx09N1bo38z2/YSnlaROAucQebMTRh3qXtZYnCFmiPG41JdYA6+fsRd
kKWa8Lz7zmR8hdTwc6de3Qk+2cmBl9eScN02O93dzBAySFwhU7/mUSUWYkLlomHceB6IdCdwGKq/MLcVhG8T/nsWMpHsXEDLK5p+JeXD5Qpru3vCPQ7BV/NJDCW0Xwom
CT7ZyYGX15Jw3TY73d3MECLgf9OzCEMljIanG/ebn2DB7Rhnq6tnp0GFIKG4dnRmWWJwhZojxuNSXWAOvn7EXVKJtvVn+CIE97RQyiu4Vlz7cqng74x7Cxf/rhzGccJ6
1iS0RRHr7ZAlYGXYL+5ly9EL2wdvNL/TOVyQyufUzA5662Ewzkt8XxXAtSVvXusOLd5DTdrSmv342gdQiFY0wQbVQoaCqpI7stQfFyd5gQqjbD4T6A6kN/SZqbbqyQpU
iYI1RWqT4bbdhd6bSfo7VtxcKQe+u2kNBhz/PtOLPtqtgMQDeEn/Dd4453bE8p4Xf9vIjME1ap2eq5OopsgIPEDWVHY12L3aOi/sS0V2MFireQsq5WbrBTCz7F8RYlzk
i/QnOz8gxOJ6k4GYw8j+kIQ+ac2JI1VCjd/9nEcZJgQP/cY6+YI4Ot88uxj5IUQylzAg3NuTojdT4wGlMX3Dm8sLguIuRFgOH1ziSro0av6JgjVFapPhtt2F3ptJ+jtW
Gl3rYtXhb5gnMCWuttfd5HmBZEzoC7CHtD+M0m9JskMd5FNZZ5SrVTA93mGsJyB/3md/GfD5TXBVSUpWGEOQIun4reAut++1TrttGg8HhC9E29D3JHGskxIUD2MWuBHw
3ZxRf6QF3YOhXQCMrdR0vVtkL9YY7f821WGSpA0Ei9/5kfUZWeGYJUU2HJ5oU449nfiFyhfjpFTD+KwxuzNk7Vspi2PiLJWB6+CZgZxH7LNjQyQXC0//OH4/kollExXh
bypdxhkgsyW9VATf+QdqOZcwINzbk6I3U+MBpTF9w5tXEFxkBVw1rVFLsKW4yOPERfPmxAmoE73AGyF3ycTES7CN0IbFPQ2shgB2HKfOl9dTp0l2JZva1haZK6GeLdmZ
KbHKa8q+RAeo+AYnr341FAldUVrs+m1751TMVYvoJ0KepePdD/AWsAFgsb5l7KJaegq+Z1uC2df6Ghl5tDjk0aE8UG7vih2pL8NrtBdIz7Ifuqyez7d2uhs6v7M6pAhb
L4kku3LgX6C9i12/bkUaMgxho2El/5iYVGXTBT8GY9bmQ5eYWCj7qkTYrVBGbjIDGdL+WXr3f1Bb7g/mri1Jdk0B9gFpVrstwDG21hp63+9KARC5IE2EUykJY0YlHwKF
mO+ouxTamdaZQyTs59MV5IJ25f5Bw+Lu1bVQPXIVI8R2ys9Cr9zonVd0RnhLqdOb0X6uGZ0VKvDLij+VoRX5YENmpPEnd5c0E9pi1kDmTljjPVL+5DpNnkkgTUz9bazQ
gL2TugYKwZjafjeVOcVBdf/UdDZLtERxA4oMQFOxGvKCduX+QcPi7tW1UD1yFSPE/7PfFfpI7Dh7A9ym/f89UfYv75k6c19lSEP1JWoeqBniiwzxxXAYtT8snuuE1GtL
Gi/c9zzV/IR7rWcN+dct7sAV8TEKz//tCebvTQYOPIq+odm1fR3q72ZoQCt+yyzaFIRGTR1d+ruiLfMIS0xOAogHZbpT2QiAm+Jy/830KVgwPfsfUTxxVSBR6/ximgrf
2/kCIcUfW+/KLSRTCF06YyM+VMlz5oTs9LOu6rO0XGZtbDoXA7jFpBezjXwVXHJDiXdg1yqnV1/DqXmuBBeHrhTS0Uk+x5fKCSUS6cGMPXWjyCRKeiQyfBDHyIYqHtfR
uyKulpYJSdrUqrEGevDm6v+eYzXyacrayGcaw/mwa/92Yxsd0xb+1GSLkbcemTfz0TFSnrNlkIRjjzBl88hxPckkhBc7pLeDIwHFK8lEtxEZsa9E1WnrLgqOmu0BNrIt
tr7vx6S/1BXwx+0ccaPKLTQ0Ez9ykQ+spyCrST3kQtmb4CA2V+dcQgmSf0WJfhqMtRbU0oksHgtPlsNUYbMgn673KwfiyfXBKNEcpCNBxR9A1lR2Ndi92jov7EtFdjBY
vESyJRpGqnHxbm/cCv7bgBfDLWnfRQJgQ1rw9iXU0f9lL14oNYYl8oQ4/eLCFWb4HOOR6xKkWEXa2GHLYGePp3MlxwlZ7hQ/GV8qdmFT6UyBhqd7mg7HCDDDzVzMt9mh
Q+w01OJJfKh1N5LQB6682E/51AV+q7DWlQiuFakfsv44DUzeXm8UDRERwKPld/wLO3hZ7Q1X4u4sCJKYOQJXHLhjVjEilRQsCPFNS4TArUG5bwLBDKTQOOMpl5vf5G9N
k61RoKCUAvrZevL8i7HXbSNAfE8s1V0GiHixYgZ+wB9qBR17tWQpht24Vd8GxHAh4gF/DtCLH7uTUxDt8WplwIj+41bml+OhWPwdisz+wZr/K8L54tRWCL32FHSHxPC/
5KVXc/wpOyelg6wbFq39dhB96TDzVV/N8EYyFHl0OR2n7G2L1+gBl8Fn5NwW8MjawQUkPG0K403lDJ2wxW9Xc/XLMV4xiyb2pGpXQ3cDteexemehXPIRTMBn5uD1SdqC
m3y1n2S7VqC5G6fzvh0sIFAvmKEH51EDlNiq1GNr+ZPUeGJZ8BWLCzx8K5UKVCm5sPwP1teQEugJSk6Rt1qejq2AzhoFJAVpSG6zcyZ8KULQbmB87tYx1Dl7pLP2R/W1
5IIwuodPGlFA+aLaW068ebLJ3Yi2vdIczeKx6SrLds74OOrTJV6rEojaKJ6FmIFpnD15WU/85ZHMBpTz9s9LoJz1k1phJzpIrGPEJhOK/b6P1IyUW3cHE/ApyD/OYoRP
ZCIHzwVmT8qKSNzul63FkCMJq+5O7YrKtKdhP/zilMR2uaY4znoz+LCrRi0l79Ycfcm2hG+IOPXPFN/6VeGMmWgEamL93JUfotuLWN788WGKu+t8sbYADGua3ezHvns9
ZCIHzwVmT8qKSNzul63FkCMJq+5O7YrKtKdhP/zilMQw4T/kO4wvMf4JwYF4Ur22wvgJJ7ZXPeNACHGIZ5ucLARUgGa2eEOndiU6Qf2AXRVT7YkxStVAurM/0dhlxncC
iS5W1jiqXZvBqC/LtjWzP+EVeYBtHot7eYFbO3lBiAEdRog0FeCbNMWTpt+ES/6SfPM1V+YsHyT3Dau2AgchFTIjwhvnrhe0lNXMhJVvYjtjULoFZVG2phyu+RZn9qpc
uGMMYVmYPw38oSKjtJX7tIRwugVV5qoH09dInWio5ztMSfThQgFGO37QJG8CwJeU7O2USWhCd8WFFd/0RTomK5mpe1gDXeE5jz3jUudqJD1UYYB9BtIav2jaVylkJsp5
ZRkdq6YemoKJlNjmbPErXFP0tRPzLws8Af9+qDMDjqdOvs5Jrxv9PNTpNvWv6tYEueado/qr2IQ7sDdlr/9JF9SBzINW8PDOO0iSqQaQtaliHKJpEGqUPYkPT8rL5D3W
uKcgz2ecFIVwzdewrZka9PifYfiqLxgTAmEGvzI+Tvfwz/SoJTVXc8M6IYClLu0LWAX0aSq8jdPnfYofg3WoHcTv0A+XGky0d45wttePIkAU5Ihncfw0gatvceOWHAvA
INCra0ICeLYWqYC8KRGd3k9w0qZiybDf7bbxqkOxgkEdDzvCjNT77i2NpjkAPOm8n0ffZs9+wWBCwzI0Nz6khTs+FcowHIPWZY/nMBcBQ17PzCzhiWUBIcZVeg9pdRDg
NtXnXeVzf94QRinks/40EQ66EQNR6IOjts6dbUcg9bNRovCvkF0Pm9LnK6U/f57TcohLipBsUL1t9gqJSGPO3TVgFwCgjHl7azLRiJpYD/mez9l7f83N4+GT82oLF3fI
1nY9LwffoMRPN4+vlD9guZDY9Lhzy69dyVTDWe9vyCmfx4MlcQmg+g6UHyM4v5ol9u4ieeKj+C8U65tIwFLHbPjaAJ1Pve9ebeiyPu+3eErZUBDE4PTEHpCPIxDq/qux
f4q4AGI0Wqfdk49JaC7rm2pPymAHnhPCBsSCoszBJ/UhQns3zaf8fDwA3XqAqZiv7ZAtWbCeVEI6yCqugXP3zdvlNqXOaLJaYT5jp4ywZqBEOZOp3X/8oW9qzZhNComk
M0yRJkv8JIwwz622AY82yNF9Rfk0m6jH0e8QTgjFU5Z4KRWldZIcMH31sOXYguE8dD46XOsaf67vwBMz0Ua/Z4wMZuZ43Gszf0aU0WkT+hFre8TtU+zEofcmmDhlzTFV
i5sEJDsjSGyszwCXMa1kLgUfDkhdbucSpvpGFqvJEHyVJdnyU/Dre8ETDdm/hv+bUO6ItKLGPLA5yQ8KYUPtJfifYfiqLxgTAmEGvzI+TvexX3v5/ATtDgpllwZaz4C9
DaCxRn5y2rEHEv9pMyZqi7xV9r6a7EmuVY8+GRGzi1iiKXkfcikkQCuO4VQjYDp0t71fFIgTDTU9g1tTXr6k/ai6AJOnJ80ywR0jDExlseMQ63ZJdBPsibXI91uvzeQE
c46Roo58kiShsFqV/xjfRiCyNABaZ4uDBXoVF7P3/z7Z/2iroB9WySUr31GSHQo0teVfqy8XcNixAQQ3WCAyKbGv/mPAkKOEcjKgFJFuZ5dNTnVK1C8ETjEaFSCCP1k4
/dOnc9OYw49Fhnhyq2gtsqIV+qP2bivj/7M4WQDvMprlTQB9mldjqx8tqq0rmNH7jDKIhn/JlJN0UDCgQYdezx8Bd3bzLW7gHX+IjNjickaJhc8rYq2iPSaLPU+tCBSb
INCra0ICeLYWqYC8KRGd3nMlEYz6RtEm3uQU3Ug+gRl+mGZK9qqCi/xokH6xDdf90dgOdXOCstXalYh3Q5Hvruu9iSp6hfStMsJxhHyV3tWZ1evTzjRo3Ct1sAesZU21
t769hW3afH2KLWPTw1QK79+qX1+C3d/yg0Ua/uxO/LmZ1evTzjRo3Ct1sAesZU21DvyizMYMW89FCvSZI7WWQ/Cajy6A5h0439ik3anQK7pGiMCQUvYgZGi6MXsDDK1e
M5xEem2TqK2cIC0m/9D/f2uOQEBPgr0W7RC39cz56aI0slkzNUmNdg//0ws45uCIxJgT0pNCgmeSk1QS4wGXgSwbFQ/9johIwJp3b8jlG4hVseClRk24kNSfzvWrr4pT
Y+KbJklH8X1b2jemU01fkTdm24RxZXn22iM+8LCY0LoyuX/Fzfz8Jx4Dzw/TjjBwdJuBBBvZlSde3VhOTgDmfy31XsPXBe6Mp58Efgv7wZpQ4UnBkDIrATBm7se0jqV8
FLTUoLhAhpEkEwBLF+loVDSfjM++WWV2URRVjJBZb/ef+GkfYiIalMywY3yWE+3voEdAN9b3CcNkNijPC0UnZB0PO8KM1PvuLY2mOQA86bwoK4cOJeJnz4tdPXSIJsXz
7PM6cbzV9ZpRfb72bmTG9yxJdtGiWVmD04/hbAN1AQDSTGeObs7fK9H/zE6InBQ5tTNEPpTcYh0yWk1IZlzPJzxQogrHIgddBkz/1N+H8D0wuAcpZgVhGHhjwoElgDSt
Y6NOa/iaOgVWRZQJjValjh0OcNXhW9CWE6yq21HjWOYl7YHFRa+1ICsx9FOFR1enWhEeoCF3s0/bYRQKB/YkBrUwKUQ2Dfx5jZBqAnx28XeJA5+2qXTS9YuVxbXIkN5p
4h49K08aGem0bm/AE6/r5qFES7r0Xj5RL7v38olchzAseRLfpGQB3peqK6cZXTz5UjV4+ImtmplooE699ttuQ5bnlCY3JyJkH+xrSPlVkBRM4x1hVrUC73d5DN/0niLC
GMs6hfhGtmY0RDnZlU3zNS3O/Vf75ZljuqH7gl+KLh9Lc0or+yHW6kWHksI4xOLcvc2DxPnBxd9/9l4VqLAYCK7IJwfc0o2Lng6NZiBdODkdbxdAYTi7fuWGND7U1ypy
3FLK9zSVami7wGsayMtC/lI1ePiJrZqZaKBOvfbbbkO5sdlifc9Y0wYXx+ofjcoKWHksVpJmw3xBTMD1kXi9C2aFAAXh82eNWd30G9SKiPlOARCoFECOYCIF7LXTh/17
t4tonZ/uPsgF1gg/bcH8qzAH322Rgt5d6gSX0CRXjMoLvK0vxhu/Q6YZaCc7gg+Y4BbcW4fuHBjV4mdJrP3wbMWSJn61vURAlBlCkYntx5xzIdUCK3kDHhi4rJHDvAUg
oEsThpLbA7aesdVcyxh42MqIJtEmvYeBjKtfeWMCbYi5CLEvxaKDTb/6rf35x/GJ3FLK9zSVami7wGsayMtC/s21e3uNNctjXEmUDsIaJ1aDZ63cvbZfXkCwfUipX5LB
N7iDfgqKSBZM9YO80p80fI4nh3iHDAKqpOFD8U2jkv021edd5XN/3hBGKeSz/jQRrf+gVHrDKNe8tpy0Wy3n3K7tO3Yitzc2o9eNnLwa9Wpp4YVpOKgTUuPCpccEQjj6
kN1PatxQLn6ARD8GGEf79ehZzYfcLh4RSzxUNzJccZCuyCcH3NKNi54OjWYgXTg5eqQrWXIBoAB+7NOJlFZWkwBRLM+sxVIT5eDZO3eoAIwA6XKPLH9D5UrizSCa+8e/
WURT/dqGSZXvcryYkepZHUljJIlaWr6pdZklHw/CpvTMDtF2EU/qIebuBpLkh2+dMKYMQ75ESJ2dUkY4ydE4IAZ7+2AQ1M34sHSbS/OntAOcIs4p1i5m+kp6YtcRDKgJ
JBZ1+iQkZKT6zS7Y2RjhCE9POHPGqT+Ag580CVAFrymz2aIVgUoh0i1k9+mX14VNk7oWfMxWID92VuaaiEqVRyjnynOcVgXk6jnfL/a4Trkn236d+mVGIvFd95o667vr
rKlNLMrfz007N6MiRMJf9wP7bJg+P3fICwnMHSj1qAoZI7UVv25OOtLEq+2L2vlHa9Nz1nZDtNO7R1+5oTAdjYV68pXTQKHSCE/1Q31hnHdiriXrsQK4R3D+yr4Dc9Il
Hhc8UzSwCXroboW8cpIdwVX08xnhOrIzOmhBFoXE64MBXgaIPbRvR4O9HdPeJeP/J47pl2ML0XStP03yW+n5SctwKW4WBD95q8k8KNWewMCYtM7VvhrGtfTprfzFoEvy
pbk+phidm1mtVBgM3h/92JGJbv4SjrBPWtjlq+SzwuLTb04rnH1P7mYWikSt/RKe98txsis4mjr5pO1zkgOzyupB6t3Nz35VFwf+CtaW9fk/+D5MMUYa/gBYJKGaK+MF
Xtz2fFacxULB5FejHsD+IXJw8Vj2iC04fHzP+xUom+l+m2Zay/5KlIWTJhA4CPL2QyfhrU0PeRzyoz5dxnW//XWLvpPIXsFJKHvsTb8kerNJlp3uyfSdhJQGxVnQil7I
nCLOKdYuZvpKemLXEQyoCYsQwkQOv8RzzQVC93S8MK3QxI/OvcxeazATqf2OaqbT8yybqd8f9mfsY3cspq1xBHNwpYyjVlD/G2pk21qKYZTrjTWr00tp1UUw0fcEcg0i
qYCjvkbzPcf5f4iHE26QDzhmydVyAhuMyORA9UW6sI4itpvUbcQf4+NLjIVECXGg9hKeVpE4C5xB5sxNGHepe+0zVXzVBaeAWF+Q7r4XkvUB13kdxgu44M9U0jvoW6xr
/imXFIsacn0i6epMPv9y9jZfRaVX627ZhRHGzENlmPPtM1V81QWngFhfkO6+F5L1LgkCsLwuWogdcuUjX1rPaLmx2WJ9z1jTBhfH6h+Nygra0BmXWJVPErgsGRbNXh3r
uTHwpjj53V5y/Tsii+KIBalRFYilDzJ7TInlYsiVdR6mT9Qh+NdbcV2hd6Iur6ksue2MoIo2v3bbsS1jnTEbAH4wa+9dIEx4cehVYCidpDruEaI1NQg37u2beN68uQJY
nqds/sbMo3Ugf0hViwMbZST88Ehzsa7lwbXcEsW/G41aHvYYuYQYVaRNFPoTyDmZdZK51pJnhGJBVcTiMgeeu85oR2I2K1iyzuRB6WT0RF7WdIhpDdQu8yo5cvPqR2sN
W6AMpoQBQz7qlyfBccrzCuqrlszh+AtsiIgJ1mMGVqybpIA+QJZDVtK07xG+eaesRu1eCmKECu8pK+PNz61YFcJZVUkwJaOCYLoHw9WLMMKoKiPS84Bp0VXbQbHOsujn
kYlu/hKOsE9a2OWr5LPC4oCJ2gmMi5aBYYOolsDVh1iBpbotlhXsSgF2lBJ5eEF0l9PoKBABApeu4IKd613Ok2uEnJTTl3gVs7guh9Wl5gVUnn8zoLI4AWPiZAbc0LwG
+kyp7EQ3VIGRE6hCYg3azM+tdAAMxOqh9dKaddvNhKWVZ5kyiRMkiDoAWhfgdIZpLsnuvnIK6USjU9vMSTOgT99sRoNNGp97JGIgD8nQWBo50e8KruknluWs/4OuBBSm
G6liRCwI1hkJgyJRFV69/rUiIRTo59wOy0zSFHODB4eKJuxxbA3k+MvjoCLfKzXnAGt2rhhe7HYVspRENQtRXbmlfkWALU2tEPgEeq+dPi0M+7rJPFGNHTd8SqdPTqcZ
ue2MoIo2v3bbsS1jnTEbABlFqyozm9NNE7WvdOEFC5MJIZllGsjOcN/4E9CXuoWROJ9nTqgh7j/GgO+434ge356SDEwxDIr09lJe7jyDkhk60XE58LY8TPqPln2x2OLj
Iatu+YJf0NOj5cGvoB9Sban/qIxg92OEp62YhEu29Z1MK5O8jKvzLhZ7gqcL+qNKWjHaWkoG8rP2HnUvjmjcGliiceD1mqlmZuXVVqvAHfCF6apwf6mqVQz2Q68XOyEI
c9VBuPmXnWpVgNlFUeztykj9ChsGQyqk0CAOUpIx61d91L05Q8MyJ74ZBZnoO6odS3YXFaiB2eQ4Gv+fO8pFDH4la4N/vR6rxjMrdTqC9Xngzu14vjs6A3gr+Psa/kev
SLjQLBK4VSuJ50X21lZfm2isBGO8/WMYCs2JEMZacgmJl3TeNgf/pix+I/JOPhUrEw9oshRs547tkMtiASEcG7oWIGHb1wXCTVWL+SU+4RyDjlxFygrVe6ygvSSIG+Pj
36tteGpS0tY5Yk5KnVgZDIK+rz1g6rYyGMwbzB10DTx/EnbjAB/CwAq5KJ3i2IXTcCD3YK9DduRQMhnQVgyJSbQmaNoSQOnNENj7LrS6SrGhvVglSnhPeS5oSn0GHmJ0
/AXPhhJdPHskFdYEzabODx5KlGXRhyec6Hiu0N4FTFaxet5jggK0LsS+ha2JOtj/osRY8unzhY5vICYh9/lF1tRdZtkPpb6Bb9mtQ9G5IqUgG/mhM8Tb99DlpqDduvqf
fqex+QjeGppAUKIEFScg6cspFmkH//p50IseAmS3HG6QupQ+PJVq6tIMo7MMqPrixKa2aV2le32zUOxgi6nI9wQZnVu1hDprDR7vcZUN8t3kxWl6rZrY/wCJhm6JXEGq
vBbQYNflcGmKYsFN9UEZ9FmnH66BZ4tgAUtzROEncEZgXiQxSurdJLMm+VBdpen4c6FJV8bjysmwIXI0IOVTmXa5pjjOejP4sKtGLSXv1hzT++JX1Lq9FC6HmpeRivl/
XrvRca+5jmb+cXtnErI9rTIs2vYICF4RvTQimTJK+jj5AC628O0WPXGvDjO1kvmQirvrfLG2AAxrmt3sx757PUhb3QD6cVSkK7A9zVGqqOcWteuvgGYST7wRJYw2xDG7
oUvDcTciB7VS6toBsv81aSU6TDxuWpHntdShP/PcxkgMSoWKrZWCoBSsw3rDj5NHmpr40Q5KocEI4sB08xlH/RY4pVLafdwKyH01TriLrWvFmdqj0e5VEBlfh2/6bcaU
x/209W+inXJL5K9Sqdtf0Kv1pxKuI2wIUy23H0gq7DDwSP61pjYYE2VvmiAGFO3HdbjV/KI/ydsi6lihiLDzYdJo8O/705csYQoaLWXC/mBRvB5ecLt9k/oizvFdXTgL
MaUSMO1erd+LgOvxPTNLnXq2jHqek+fokHjWWPSjMrssaRbXEiH5KrbmS1mE3N0M5rgSStT4NIeyFQ4Q55W2N+RZ41RZ47L6j9FcM1ftjKPZFJEYVKbtccWGJl2WYCTt
8oQQg2VJbq/1SfnddSq0iO8USFSHYk+j/gGpyjxbV/LA7hCs1kk326wXHcPkfukPC25uC7QA/8cuVg1JlMGkD2uOQEBPgr0W7RC39cz56aJgaGRT1fiTmilGtX99BOvC
18rLA8NGlRhz8I4/AxL3naIH56/mN+Of/D2XL9C2XPScn+R7oRdESr1gvQYj9KRcMDSD0n6RlMtU9SWlM4aG+pvYE2HnlNCT5vyDAgXs0Wn0mi+gZHkZdo3fV8ANzOGP
5yH7G10FFC1zNWcVIDN0k3BuDlgVWLQFoTFhBuLVyavjtR73Rj6D+HTGArSAtkvjYGhkU9X4k5opRrV/fQTrwmLZEhaR1plDzfRfKPADeyr6DzHvp9ppydEDUV4vSFiU
Nl1E2cuGzVOtRfFC/qy4gShjCialeFGfuGCGETt6jATir8Hw7zTH7MCaJq0jyB+GpXKHsJV0YqrkbXM/od8iOhMEN56wshbWdG5P2fnJzUi5PDrCkQxNPWnJ5/YcHnLe
ijdlabzK4MRgIN0035r7BWu+Z8LRtK1kpeatUaGlilgoYwompXhRn7hghhE7eowEIkBP+7k5MUqIrFA4vwxtlBdzdryIUDjmPnB2blSe6/UEQ/FwuI2va4bC+FuhIkfv
EjoiUTVLx9AvAHDuBtrVwLw/4/fsFyhKZLrZnhI5VtuLJ2V2PvCiEGEO+KqrUptQGCyxX/nMO8GWmBf6goTmu/ifYfiqLxgTAmEGvzI+TveCJ9a1TSHeHEXMIiVYsE49
yLVZQN/7EUHvj2i78gkCc1zu4R55P3bgtmlTrXX1nobsAF300tmjyI+L2k444QJ20HNQNbrADMVsZEyHD4jzBjnupGqaHE11+ctL5I17EHLsAF300tmjyI+L2k444QJ2
ZEkljiuTsidH93CjhXspEBCJLOS+HkbD+vejgUAUYcESJHaANvR3/LgKNPs9OH+KkiU1XyAZIKNaU4RhhF40xn3+iWyfCJwL2pzl7Io0ges4XaLbxzNx5fD3BpaHiHO1
Xoq1TQmHQiDmkgEM+viIfpcwINzbk6I3U+MBpTF9w5tRtRS0IQUSvmMRUuyP86LDIUGRawORppmboxxs3g09DtQGJQXfl7N1SoJ42fFrCv3j+ebu/uJ49LrADT3VvUVj
Fp2cZ8IVuxCWYl4C5HnFslo5atVqlH38iDZayGtY00oikT5m6fuGXpwlxz0k7t7VNKTs2nT4U0g/QjvQuANJXCJViZ4LhKL1lWTc7Y4MG69lXtoVXjVMF/kGBxkg3FiC
lzAg3NuTojdT4wGlMX3Dm+nDkz3A6YbQWIqIHDSbQBDR37qdzHA/b9I3x6f/Xfm+P9qrET6eF7PH4vosV2V1J92cUX+kBd2DoV0AjK3UdL0QiSzkvh5Gw/r3o4FAFGHB
I6hXTUvv6KBrCduTj7NNhteE359epzsGva3IPotuWzc7PhXKMByD1mWP5zAXAUNe0YFeHtsYByd6s/YCfGNrrpBU14sK81Vyz54tGhCAuDzNzqr26LBZADP7KUNUK0Wy
MkhcIVO/5lElFmJC5aJh3CTwqz35Rfvo0DTcHDs0OEIiMTUZoH5Ce83m3/DuwrzKIuB/07MIQyWMhqcb95ufYDJtoNHfw7qMFs133Qtl1vNj4psmSUfxfVvaN6ZTTV+R
xD4dj6qtCVf/oHiMMOjruOch+xtdBRQtczVnFSAzdJO6hPYq7O50UYdAChllknr31eLC6Jvhtty7WJfRMxP+ZI+0Vtpv8t2IsvUSYmFHGmGP5vgk8itbiF1FMhbnHJie
boqsmUeHNtLEj4PX9DZ93sV2Wj6W8rtEDX0T97ZG8RRE29D3JHGskxIUD2MWuBHw6OTVdnE2FyDiiztZEhE9ulDhScGQMisBMGbux7SOpXz5PbD0RDaxZu7+XkzhLnoE
Cjqe27PCcvUhNrC7eXBOhkxiSNMQl2C7y7UnNBJ54QgM7gE7AGYFG4Yb8pAFf2Dmj7RW2m/y3Yiy9RJiYUcaYRsRbg+GAwLq/HFndivTi2LABW2zIfu4BoHD3Ea4l8kz
MiMvU5T8ts7YHaviRNyHV3Fa/2wetEa233/PD2aFmRdXE3UUzBFTw/0Ehr9cC55ddJuBBBvZlSde3VhOTgDmf7JyTZTxAWplTPvR7xcfYOyb2BNh55TQk+b8gwIF7NFp
upc14gCvPCyR8F0ms7E/jW7EZZTwwWo5Py1cNVOIyA/j2KSvYoMebAYY6iiN7r3P7bDVI/UqCISbo1PN3JDmto9njZONUhFjIknnBWykUzkJm8zxMW4UKQIE0Yv0qo8g
xRHvM0Vw3FMAfF+h/if/+8O97bh38i4L6JIDznhegHsypmaq2Ac+xMmlIMFLBO4NBvPbrUwtcUxCAToS9bexRLKeu84qTO2WaulIMF/wHYCmw5iqvzxG4vpeLHoN1Ek5
LhumefW84YAiQlXszupmMAoGwkM1er/PgcW6/yWpSs48jHbvphj6pThPAeAaCkYyVm9OkvSOsbbkwxZ3UT/H057vSXniLe69mVBGAmZASRD4njDMv+Fx9ewr7PfXSi0u
7dryamWkn/eRdup4R2hyJINkFkDepK8FmJUkuUkhBcgGP1nuX/ipaAnALrpnWhOwTwe2nsdR9zOcNiVnLOf6tOwAXfTS2aPIj4vaTjjhAnajAiC3ak+Kq+HeMitTipUd
pAsKyto4BNuZ90Pph4PU8xwpACG5YtG38HqqHpXEnXmXMCDc25OiN1PjAaUxfcObBfgd/TqnXZvQ21fZNqbayuch+xtdBRQtczVnFSAzdJMGJwAmnLt895XVsDUje9pT
1AYlBd+Xs3VKgnjZ8WsK/bGR25uA4DJ+DIjFkLkytMXs5D9WKBVMdqrsenEcMfBhoRD71yvPU7mvtU6oImrYYQRGL2R7eXxQSGKxZmrYbmntC2jidYycQaEjacfnw8oE
3BYAA3Nu0BMXtZ60286uGpHlfUa9zT+LL6BR9WdDv6xi2RIWkdaZQ830XyjwA3sqTmN+0YDXAjasm3Gs8MEHj5VYURojG2peArvAJeQcrWyW47nuW8c5snn9/qXb7YYf
b1EWY8eP0jWzHqug31zpWGc4pa72nWUGQh7HH2zGPRgqVu+gE81FRlfgVw4MmR7w5yH7G10FFC1zNWcVIDN0k4OFumER5ifeU6o7OgQFeo7nIfsbXQUULXM1ZxUgM3ST
h5FJWXqnOJh546AevvZaKuwAXfTS2aPIj4vaTjjhAnYV7lic2/rKBTntqlt5iER21xQpONtnWsNvijx5cvFdwHLD61xHv+ffRNZQxfXwHjMqVu+gE81FRlfgVw4MmR7w
5yH7G10FFC1zNWcVIDN0k50YUHR+TWRfmgzv4kGKoOMoYwompXhRn7hghhE7eowEPPA25TUymcMBpmZ1eEtPmu+8V/DsAatiYXlux28s/N6Nv1UY1/6OE20pDi61FOaw
hTSCBk9c6u5IyXhfNC+TYSM+VMlz5oTs9LOu6rO0XGbskI+DmlpY9zN6y4XRLLMk1xQpONtnWsNvijx5cvFdwPnsi1AQSeYJUw+lAFQPMddE29D3JHGskxIUD2MWuBHw
Om8btGrUEib74kKFF0KlM5HlfUa9zT+LL6BR9WdDv6zJkTx38zJquLieRZiUlINhEbdxfTKy4max+WUrLne6i7ubORLeiDWDVQfwFIsRd8R+Ag0NURNi8ehVA+0LePXh
d+/ltRNHyDKKFjMp6SnyssHtGGerq2enQYUgobh2dGYBYpUlBInpWpnJxKzzpAK+Uom29Wf4IgT3tFDKK7hWXFq3u/7iMS9hh+auJDVAr6yqGRk2NKE56JSKxKf4ePQa
I4qrWzg9D903EzYqbeuSHxsrlKlVBtiWM6JWcRhUHOrcXCkHvrtpDQYc/z7Tiz7aZpVM+5OsccqDcGsxoFDShFKJtvVn+CIE97RQyiu4VlwjEw6Rs1o2V53wJxSf8lhA
ooelsXGfLkOi9pPYGauRLOGyB4FFotbluXPSe/r51qiR5X1Gvc0/iy+gUfVnQ7+s2/kCIcUfW+/KLSRTCF06YyM+VMlz5oTs9LOu6rO0XGbRC9sHbzS/0zlckMrn1MwO
I4wTvthVF+ATr5q/pKNo5tkEJWv1V8aH8oY9VMasQz3NtgQn8+PHOVhl/FMECYOUooelsXGfLkOi9pPYGauRLGC97zKY2QP3jtmg5o7+vAUt/U+a/F7YSOjG9tC+VAfJ
XSXp2wQTo4YL3abHgmtqK/4uWP/FYdWLqwFDU5osxVeiX1vgGnK+6RkNEDk7n1cr2H0MSaZ/xLBaCHRkHT6AsPXKUcBr3M1BDnhoyplDtN5nxdgNYKcurSLoAg4DdLLC
kTYUCo8ne2MwD4wP/SXwMYX4yNemh6dyy7Au/izbrO1NvEm5+5xiXK659LkdGWoeX9CQNcqVuESgiK3UwmK+um7E437HC1wXcmFcnlY+Hx92RpBI+6WK+Otjit3vABq3
n4Gt8+8X7V2RYSIQ3e2IZ1ePFD58rCXxIwo42G+BEkYZ0LfSgclURtIvtyFwQLu+me/vEMZY84PTR6Gzq8u44Lpwe8lN6OKEQXleE9lxcQcPs6/cgFfUz7H7QYKUqud3
uTd2mmaSU+HqbQtlBZznX8j0Zx/EVFFlOopE4AUtzhXsRc4a7+Py8x6d94jcATRO0TK+oFXT0uDCZ5zvVimHvtL1ByUrUbj15S39JAdzuAbN2zbtICS7LPpyY3GIS8JX
lShWgJzQUbnO5j2K35n2mOhM4DX1EZIqEIT/2bGNPdwy8i+Uo1N9hgwDrR0VUglwG/g/l5g1iyaDAlt5dy7BoLXrqYmYYDHglc9iTY8LWJbNbfaOspT3Kj0hrA5RDCuc
Q9GkTbX1FmqJKnY7kPwUoGuOQEBPgr0W7RC39cz56aKYUSCjMmGTYf5Z2prfc5i7lmTBv/Jsyh2wrXC7dMiOos3OqvbosFkAM/spQ1QrRbK9b6D41irYa+jPP7O7E53N
hb7NBUMJAj5WnkvUVcUuPUMq+fSCuDMGwAbQLVTLjMLfR0qMaTxAhw7xanPcz1Bh3rR8GBKbDIJp+vN+9qM9lTxfTxpDPkOaPOET0WTILuO+griuZYzFP/q5+O8qdiFO
frh0T/LImH+xiQ9SZ0u8Faej1zBicYLRTygtrh2byv5LFlgBByx074BnXrQQl6mlAUF/OzXG+4CG6sl050Lgv5vYE2HnlNCT5vyDAgXs0WmxTSv3+brr6Qqu6Q3AoPsa
9eOACL92mWw9SMPNnjPoCXbZsH84QoXIUoelJaVXQQ6YrFstNwLjW6zaf42P8Q9QYx1WpJG7WD/Ii6RtrJWMeCIxNRmgfkJ7zebf8O7CvMq3MTGMZjn3Jb77jzm2Hvnx
kuuhhq4mVW1kDGh6tUBNx94I8ubpKt7IJYSwUTeG3LzsPWc6/H8A4yZuiW9/UlKi3rR8GBKbDIJp+vN+9qM9lRX3i+4Wb0MOtHWeSvwCSalIBEL7VufQBhr4V558HR73
HHFmLwr4eHi8nGNaFJfXE44p/tMCZI56aY86Si4UYzUuYpGIjaUi7tf3s84xauPr3Iy6qz8HQS/7uDhbJ568p1DhScGQMisBMGbux7SOpXx552et238vJqaJkbGMsJgF
OhO3FOkyy1S0YiLmRltveOO1HvdGPoP4dMYCtIC2S+N4TU963dWEzm5+3kR3EDBnWAX0aSq8jdPnfYofg3WoHa9EJowp9vyrbrJHo1fMBR/a71uD2T+u15pW7xPs3hAC
a45AQE+CvRbtELf1zPnpoivbf4yMoVOC7Ewo4YlBksAQiSzkvh5Gw/r3o4FAFGHBI6hXTUvv6KBrCduTj7NNhowmdl2Dz03ae5WmJvjAsd47PhXKMByD1mWP5zAXAUNe
D1n8akpRY/BpdeDD80rIWpBU14sK81Vyz54tGhCAuDxrvmfC0bStZKXmrVGhpYpYMgujrgUWqytO1Y8KZiKPoRCJLOS+HkbD+vejgUAUYcHiyN43iNeFvHBlmcUGHUm+
XNshusuSYPwX/ctHbby4hhCJLOS+HkbD+vejgUAUYcEjqFdNS+/ooGsJ25OPs02GVVpjiPqkba0cSCinAC5pwtkUkRhUpu1xxYYmXZZgJO2vK/wOLI6zs9Xe6upD8jMK
xu8VgRFg12TUBU2iWQOv6YJXpGJrU1ZY+t6574RPaS26Yr8CFjOM31i1LBJmWv85c/OShjgnYDBnHLjISR2qkYF+GUsnBAH8lKneVB/P/l1ubqpLd5nc69CK2aqexGOu
HFnRz2MQdfLjJI9RJoIdhRXK1gVVnKUAtaWNRUqhH2W4BJXQ70QUa0+puF/S4lglKTEwZGDXGFJDW8GRGWNy+Yk9S9iRlNT2wIrb3ghaNXsB+BcTpMT/2QP1vMzPoD22
SwfcCSA9Xp7cn0aPBQiRVBCJLOS+HkbD+vejgUAUYcHiyN43iNeFvHBlmcUGHUm+DL50TtcbJYDipTV5QeQ/p5Gb/XjYf1EkRnn4FO2WZFpB2DWxvY+ovEfhuJrpMvAa
ln1o+ySC0gNmnM7SLHWdEetrHVCQRpp8CAK4u893V2PMfgshykhMvrOqs4gh7IEAc/OShjgnYDBnHLjISR2qkYF+GUsnBAH8lKneVB/P/l0TxeqMD/4P3DC2OnCNAWiP
s8Gwcia+HHVaETifssqJGYE7XAGJcubqAdzL6zJAGN1Ppn9l5Aw4aC52FIsRpNYKGAAhuM2Ni9ofyDfTayGPLpWzKMSD74BZQD253+9GDdIdDzvCjNT77i2NpjkAPOm8
1P2By2dH9ZJxehJZ35mR+BCJLOS+HkbD+vejgUAUYcFnYPr6j2cL0MtwVd7kbI7afIS1wJ9i4C9LQN2/vQ3Xv7z8MYDGRqjjMivYGuJ1H2qbC0TvyNgNfJdjyu9hwmZY
EIks5L4eRsP696OBQBRhwSOoV01L7+igawnbk4+zTYZ+CcteOJ7w7hbpGO2wCoXTa45AQE+CvRbtELf1zPnpog0EXR8NGdvoUFm95siUPfrpDwEEZvyPjqh4KSNVbSCo
kJe0dRu9ydSsdAOeehmyjt4cAAHQbgDoDRqZi8awdC+oD3kUooogUi6zTOi/6Cb2zc7yhnNJOfsrctl3fb26abBn0DsEqNvyb6c5z2bmzip22bB/OEKFyFKHpSWlV0EO
If26DnAuM7eeCJagBZtjkCdUyja7QPKBfEIkEGhOw65rjkBAT4K9Fu0Qt/XM+emiLcv0iLj7hyP4gv0Y677jrvifYfiqLxgTAmEGvzI+TvexhZBryajCigs52Iqycm3+
rjJvK67JGXLZhVCwdaIEfM3bNu0gJLss+nJjcYhLwlcRlmykzWxUmoGdDb054UgaiktdMBoRdjinx5uNqpFTBN7YN+iWSI0zfA+1UPUf1bKQL042ZKgHMWS2e796lxG2
QMxNkWuDxEAUlFeF+aSP4q2WPl3UpB+JWOqJkkljU1dweAzGRO6yOaOLP60W6Md1ONGzG0Q6RgKMYNvsVn6qKuP9uRzUEnHTeJuWizEiQUylgd/ns1d6GvIejMzwtSOe
Yvczp9z2nBtW4MVJoG1QYd4gceAKlvAA/ptZU9DJnXuwz6ws4LfIaOjE8aAGj72J3gjy5ukq3sglhLBRN4bcvOlztf2KaQyxonKlOtveizvIQhzwoXrJVzFDLpHKwr5n
3rR8GBKbDIJp+vN+9qM9ldgxKvyaoYEwPzhNQOE/q+zsAF300tmjyI+L2k444QJ2jkHTfu1FqskX+HGXFRYegjNv3tUF7Lk18y4HTUBrwiO7dBXlcGF3wxwpeJZ7uJOM
oXXvS3wxDP4SYbI++QUVxmnUB3va2TbwVX3jZZnbFp4hoYLzsBKAHDg8GFjNFAvxjs/8VKtLttaKsRkts+b9uX1yEn0f0k4eSQXjzD6WjIMg4bhbVoVNR8l5+tmh9qcW
cHgMxkTusjmjiz+tFujHdRto1TruR4eZ1tECV23cD24wZW9LE5NXSYtVEf6/wNbI0kxnjm7O3yvR/8xOiJwUOZAvTjZkqAcxZLZ7v3qXEbaClkFLM0oE1dytpYYlE50n
ZrfoB95lGQNZ0lLDO2XunOtrHVCQRpp8CAK4u893V2O7dBXlcGF3wxwpeJZ7uJOM4g3GhXDWW6dgddRYU5141FXTlC8iCZEd/ZoeIRZe086vRCaMKfb8q26yR6NXzAUf
CcXpb2GRrFO7e/wF0kXR4S+6NXPrsS9R1t5kboLMOhabPHvIjiIERCJI1GH5BP573gjy5ukq3sglhLBRN4bcvOlztf2KaQyxonKlOtveiztgCEMcCJgW710n1wLjD9ys
3tg36JZIjTN8D7VQ9R/VspAvTjZkqAcxZLZ7v3qXEbYZal5LrqH2dymms+z09+nVhN4LSGBgzYA3AaqvHjYDI0Mq+fSCuDMGwAbQLVTLjMIrHOuN78XnBTUn0bW9m91f
NfxZbG1tm+kgoy6xdGBY+QoMtDSpAI2i9S57Ej8nIHnOcaF+s8oaf6ok5afGT1x5ehxJh26eG0iu/A7AE000wIAYdPsQSNKa6kThnGw14jxrvmfC0bStZKXmrVGhpYpY
M45djlhp77QHgApCsFIShA2CXiIS4PhViz1nyDTolYoA9yhQhu59m1d87351rsN2oMCTDUeHrEU7FM3Ln3Y8CwnF6W9hkaxTu3v8BdJF0eEL5q1xh9K4MtAn1HWuLvd1
mzx7yI4iBEQiSNRh+QT+e94I8ubpKt7IJYSwUTeG3LzfVQ/eH5L48k6uUqN1fvPbNplpTDK4lIBf6rIUe9FOVbscyheMGBf297+1s5w5SCOQL042ZKgHMWS2e796lxG2
RtAKUYywneD4GhcxG0zV7hDEtRqratSiZ3EM1JgNUo3R37qdzHA/b9I3x6f/Xfm+zFyB9sh7GbmpWwlpDhvfLUTb0PckcayTEhQPYxa4EfCnqVHzvrJv5B/sgErAnBd4
r0QmjCn2/KtuskejV8wFHwnF6W9hkaxTu3v8BdJF0eEaApuqJpmmJ1wxYXybaXTcTJO2jrOfAJAEu8OA+wNJcxxxZi8K+Hh4vJxjWhSX1xMCiQsqoD2HA2mvvEWfZywJ
1D3ykz9mrBRmRcH7cLSu1x0OcNXhW9CWE6yq21HjWObOcaF+s8oaf6ok5afGT1x5ehxJh26eG0iu/A7AE000wDqYeOx7TZRKpzet8y6oP3Tj2KSvYoMebAYY6iiN7r3P
BGGD0hmLNEUxIZS4DR70hyYjy7ndGF9XrX/ghmHnszatlj5d1KQfiVjqiZJJY1NXyoYCt4HZsfLXwLp7jso1GcwH71xp2I6eRNDSVOhy8XpjtrHTmPYhK4OUTFN5aF7W
RoDALxAL7WnR4RNaeUVDqpDdT2rcUC5+gEQ/BhhH+/UYX5ia1JmhOs6Nm3zgrx4Qyogm0Sa9h4GMq195YwJtiPNcoVtfU+2TSgmVMtMcuEjN2zbtICS7LPpyY3GIS8JX
QxvBWLbE6DcPmWR9oJFq3PeubT1NY+WcbifVjzBD2A9HbE8R0jHvFGkRAPbPyPGB1WEmeAUXYLQzop1wC4jAEswH71xp2I6eRNDSVOhy8Xq2b9nN+WWs/Lyg4VUdTcGx
zds27SAkuyz6cmNxiEvCV1+W9b468IDBHET0740BOnyZ3MlPzTEqdpRhzd0apuj2R2xPEdIx7xRpEQD2z8jxgfqJjSXcE9Js+zYiKU6nw33MB+9cadiOnkTQ0lTocvF6
S8FXe2+h00EgOYcDsSasjM3bNu0gJLss+nJjcYhLwlcdSOA8Waq8SxDnzh76k8/M6DVHPbY7uiNyKx6dR5Q3jUdsTxHSMe8UaREA9s/I8YEm1sMlwOWDLgMkJNf8RPM4
zAfvXGnYjp5E0NJU6HLxeoFQ/yceo/pkA7ZUuHJLsxhb4RYEzYrEFXQ7AtHw5vPl515DVbVtMTuuV4v74ry+kBtJ0y6uebPTZJSjMfQ+ZotC2SZ8RS0ftOftsC5mfZf7
TgSKn20ZL8XxbTGr10VMAF+kePubDXEHzogHEF9PZff23vDNphlbhts8zt3nTelShyTD8zaQha3BpHU1RMDmySGLB1zzL8IC13BaVDGOGVOWAXe58Nnik6REX7xWcvpb
KFRyCjG0vmqbFWeswnv7pqb4Tti+yzOWq0kjxbckbl+YfmRLux2QJB0IDHVlzi6vcgYyKnXcGPnun5d6d0mNez+5VldoF4L6/t5ZiD7tnK6SRT/YSvMWBHsllRHKE8TU
SAFok0Cm+dUH3WrtF09S6iO5c24CEo9fOl0TtLIhRI4ZlHbG5vV3Wxz2y7q1Zc9tvd0uRDyoFG95YHQ7UgVa/2AJeakVCnLsdGc1ELLzFz6s42YEf2Ox//3M67ZnYneR
bBAKYYZoMuVDposw4NVYQ5nvwwZQVl3azywKtMECyzhXDH4OzChLhvbqmLXvhM1Dl9mufuBMw/et7mXOf9ypVGiKiJ81BI7UskWOR8vPOG/KiCbRJr2HgYyrX3ljAm2I
pXDKFKryJCC7lxqSMgT5fjbV513lc3/eEEYp5LP+NBFlrzAuGvuPbU51bvvesJ8KqMazfNXUNdk5v7+qeiv1qLOBDEX0oabzdSDF0rrZf2DbvgMINEPwcf7e/tubne8P
CCSj3W8m+jzlpHQId7TLW0728kUeZ7sin9oWLIVFvlOqJ0iLlGE6LIT4mnZjzs23qOgCuEUnICXcB4NG9FH4IR4eIS8iVTQ6l0vbM3PWy1mHXjnxAIX5AgoWYncfKqfm
ZSYd5uY2EVwi9xffUXZSMJE2489efz4PPQVNaHOJFlp/MAUzUzSmBRwdz4AhLJ4143CWhqmHb45TqHfbJtTaCDWlcsUoVh5Wia7H2+g9FA9gEVAWc0377dkRbYrFLTwf
XM3JN1dksL/FmuaWh44qdXM8Ej+8WDn/41DgujYjpa2VF/CB4e11kXAINC68FMwY1NXH1nFoSDZzzJzV9cCZpO5tosKkGPxWTInUzwFmzwZ9jjpMtpJK1zNCMUbQsfhT
1HhiWfAViws8fCuVClQpuWduL8EirGTbg4W5F5iX5OmD/keldeh22oeuS0byJcV/hk2CkMhi1567n9l9qgDTgLcMjcbtl5CzihPuWpysojgqcrCYwA6u3uShQpO0NtsQ
vSpdm4PpNIhNquCWbFco0oerXbWI0C6h3No9eIoQLugxgB5OKZ4euSU0qKJ2+2d/KdCzIkhhsuF0AJPrg3eeP5onViSkwB1teQDAsSGFyzopWcP/XiVQ00nl/j8ZwbwF
HHwtbI0TlMB0NK5jb5wubBayWE9NGIn2JVQuOVOQLHnRvnYxnz2vYml0crQKQ5hK/rpTUW6FzVb7uq2Mk2ms4XYKV129+3VLTSzn8H1IaXYp0LMiSGGy4XQAk+uDd54/
R0Xtcu9+mHLOe6ar26k7kXwvSa89afTi5aYsJLmSHGvdBJGSNc9BFuaZ6RGjjG7TPIs6zofvnH1JIOBuJTij88PnQJUdNGs43FiOCb9Klou6oLUwIhiHCemEtceaXXkC
wapJFD4lnaMwtld0cbJ8Z5OizflI0mg9XKCo50kTh5KYPtIbcXosCyDXA0N4iWYDBekN9ToY5WRth/bI3CzVjbcMjcbtl5CzihPuWpysojigVJfBZIkdIPbMdMQEqT6N
7FHKZ7n9WVbYvWAn4RnzUDGSUC/FziiXZzq1UABxrxAztLU2LawqywRo0EgIGbzjJrt2xXNZ8eNufrlYiFxgVP5cOd+vPQj6E7VN3s76sjcGfgyve0lZel4iDnOC4qc2
KdCzIkhhsuF0AJPrg3eeP5GyA/4uKeXxqUzKbbJIq0p/4QeP5cOmPiEPCwItwyWKtwyNxu2XkLOKE+5anKyiOBYPUbwa0ZT45aUZHaYYzmWx6ZPnpHLHM7kE9SdNIBEN
IabEGCI08ySm7rJCQDGLiIgZ5fQD1jgNS6v4l3FD0BEh07YZ4GQSznhX6GNwYsbqG7k4cJ/PqKkIx76xTRyDBZ6/GSGYVHJXKeVQ/pJ+YR7d3dy44Sf9AlAus4gL54I/
MSgZMeBozshcFMt3ZcFOoUge4SKhEmpzJmQ1u9mLxYtQYzlQUPWL/KQLCdEjTx5yMRXwZa9NxymmiG27c2UpDaE9EN3vBfVjK+mLoSJWtYC3wXYuHLGSOx90DchZm90g
EmnrXSHPvINs6abypwI+xh6jZTUF9indFQ8nKgKjXYANeC37Cz/GYfpvcrdrzXy8Cf6EPdBfjiXIp20K3BK/8NbHSNycW3ZL4F9eoPJ5dPKvgfuqCws4CFxjTzHxNAes
S5OHQexaS208Vt4GT4BXMoy0/IN9lpY5mJY8aU85gL1mtn9vsiIKpCkKXZMuuvE5PtKUyDLjpwhqXQkWpZ0O/5g3J7u7ysg2H8pNbITOdZCf8CzM/I6g+AnFVM1xmCHl
EiRmyFlI7fWVrvsEk7Z1Fjq+zxDhT5xSTufxyJSpR8puTn+aVgREFQoWqdUOvLdv3fdyYNKT1Io2V6H63wgKobhRfnuk1a7KAvNsm2apf/CWwBZESJRE7pIecjNnGu+7
yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUZ1AB+02V5BXdjMlgfKRVsHMuHGaFiqC0Va40HOdhiyS2AvNpn3pPX6TaigvZdE28L8bUaFrrUWrJ3C8NEGi0zH
2IxgPx4X0/eBdEw8eySRiEDJqrCQCDOrgCkmTBNGpAyuLUiaGSbRvMiO2Y5sCASNAiINzVxRhiIGSrTN6PWs1gr0S+U0Xeyz0pZAxMjivBaWYnCpLHNzGAC4XS62ftEe
9eAhsbYpcvuVPp86ImPIqn19gEBZcosw71mff8zTfJfpOQwmyrJONThm8bNO2FtiKtHHUmYJBzO9SUDZlVA8xJbwzClTy4XZndapCNNU+PPeBEehDRu5tBQw9W4ARUw6
3A/HQUAYHGYwc9euKnMf/O+Th44/BTRBMoPlJd1MJT/FgieKj3bLeSCOFOyV8tz50Z3EwuRSCPStXyUSkU6wGcqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFz
nJ/ke6EXREq9YL0GI/SkXGwRJGuzlB+/3aTi2zR/MO3l2Q/Pajdjxho+bZn1KNVRVMaUMndBwF+kwMksXvheRp5DxCzEkASNymFUZ4DxMUYTiY/nIHLUaG7nhQ7jQlgh
sjuddenln8ac5VYKnkY8n2g4AHzQnOoyTHIa4yTMT+ZXavGLJ6DWVSg7vYWTRSGBT0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCC+nMFcJRniBj9+MV4li88z
cguOlyTEP3LaPcSElVlWBIvwrK+x/56RzS7EEaSPliTKiCbRJr2HgYyrX3ljAm2IdEMpVk0/iVLB/Xc8gKO+AyQJUjdB8uRmWExm8WrFdwHUsLylijY3gkKh/X990ZjI
DJQXNYxUUZgjoAXhf63258qIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0i70HRoP7GfTHaJ0xeliBg2Wy3NTGmkLbbDnI2+3pIrbfGcBtsnHjiIIwKQy0GG02E
MKS9qjr8DhbiP98e3EH+StMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o3ea9yDxSSJF3wt1QQcMeY/UOzgVhr2GoovWyiZv7yBxqqYR2RT8o3jIzS01USl5r
yogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh1E7oBqgUkTyQDTN8Kl7aOO8EdSPUz4/+iCZhpsB7CeF/nEks68gsjMbQlHTAdrX/RuPcqjj4KMfzKD264bGZmd
gRrInBgZD19HN9j5BZzno87kdbcVAiUyz7ljCbFNI5CflEwYHZwQwKKuv2jqpVYOmozKuqkViTWKEFs0tWudcFNsBzzkmI8VT8mzzaEM84/eBEehDRu5tBQw9W4ARUw6
K09CAaC+GdPoTocIAxv5eBzy/vYxc5wDFeFO2pzsq1pnE9PRDtnwCVnPJi7Ue/W6jb7vBTZr/jGplhPCrz44S8qIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFG
qJI7YEbeIAYkNBFAqjXCBKH7e6XgzvuduYi+LZn7u0II+QhPVUEsLCCU9Y9+S2JGTNaw+g53QpRJfxKWC0Pwy+cDINPdkN0IRxIRWcP/qasSRqiVp9bf6hq6IpjBQBhW
Sly4z0Sxtnw0VPtn4NIa2mCAoeqsGCXzyB72PGVSnGoJxelvYZGsU7t7/AXSRdHhkQvSanyvBAlBVbKh6MPoQut48B4+Bk09Fg9hYF35DqKokjtgRt4gBiQ0EUCqNcIE
ay7DS6XVXYcYFc2rT2jwswj5CE9VQSwsIJT1j35LYkZM1rD6DndClEl/EpYLQ/DLIM/AlvMnyp7b1++Eh9RfUxJGqJWn1t/qGroimMFAGFahde9LfDEM/hJhsj75BRXG
sbuM5xjuyd3myH3AOqOAiQnF6W9hkaxTu3v8BdJF0eGf8wPvZVcs+0N3jEMPJq02vIUBs7AlkTdVO5sdbY17dqiSO2BG3iAGJDQRQKo1wgR/lodsBscqqdPAbQkXGQyo
CPkIT1VBLCwglPWPfktiRkzWsPoOd0KUSX8SlgtD8MvQZueJC7GqmVyxhdkNqLPcEkaolafW3+oauiKYwUAYVpzJPIvrIemSLOsF+r17NbpUoCwFEL7owHPR9y+0MRct
CcXpb2GRrFO7e/wF0kXR4aB1uDZqewDNWmSw1fc/jo8i0ZW9YE28/xo0lLYLkHpYqJI7YEbeIAYkNBFAqjXCBBF1bUcFb7IWO/p955pUqLEI+QhPVUEsLCCU9Y9+S2JG
TNaw+g53QpRJfxKWC0Pwywng564rQ9UHYyCLSeSZBhESRqiVp9bf6hq6IpjBQBhW4g3GhXDWW6dgddRYU5141AiqVzqYDVqOCASAYMPHNt0JxelvYZGsU7t7/AXSRdHh
71dCMIWBe1z6ZQYcPSesmhpfTP+ipNTNECc+nUgZh1+okjtgRt4gBiQ0EUCqNcIEwCPxXrQRguqcT1WD1pk7gQj5CE9VQSwsIJT1j35LYkZM1rD6DndClEl/EpYLQ/DL
LEG9tkZz7ih0UOnVipii7xJGqJWn1t/qGroimMFAGFbxgo6S2FjIiZAxtGi+DwOZgiErpBjMSd8XR6j8KvZWDQnF6W9hkaxTu3v8BdJF0eHEpMLlU3HvGi8vEgZaR8k+
zaH4aZqWliI6V5x73u2dS8LAA8SMJD4sHLNJVt6Ew7+LYGtvY/Vs1h2pytLRB97ECPkIT1VBLCwglPWPfktiRq2Jsefd6Qwy3BTLGnHfQcpNf3RUCPmzaE3QNwrVymL0
EkaolafW3+oauiKYwUAYVtxvP2XNaKMs6Ppux8JBg7cHvi9svv2sIBtIX3uxjDSAyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjTIZGc9kTWzrYMDyDvnYgc
uc/k+OXiweAW5ELnA4Vm4MljTIfYsCq6sEaHJiunc2e4YWjxaqk39rqDGQqHunr9Kxzrje/F5wU1J9G1vZvdX1TsZmG/xjlD8L/OUTqK0i2JC7IMZSw1YTfxa19ZyEOu
1VJ5bDR1uK10cJGMv8Jio5Fe3SGfe+t89Oc4F/fdbLTMXIH2yHsZualbCWkOG98tRNvQ9yRxrJMSFA9jFrgR8D/+yQWpzwVNklE3mIVLoFOSNw09cGng8UC0zuarcnzV
EsSzcNPaHZ3v3QbrniXWr05cCJ8GOs3J68V2MGuRpUsrHOuN78XnBTUn0bW9m91fFNhrSGCVVpYL3ESqjM55yJcxlX9YO+c3TxxC0LDHZG7VUnlsNHW4rXRwkYy/wmKj
89CR5KVNEaw9KqOqIkmdMMxcgfbIexm5qVsJaQ4b3y1E29D3JHGskxIUD2MWuBHwatsRNq43z+TIsPBtCPExRZI3DT1waeDxQLTO5qtyfNVKtdon1fV06N8NgVamJdxf
uGFo8WqpN/a6gxkKh7p6/Ssc643vxecFNSfRtb2b3V8XRKkxIPoqpes/yrAnvj6ApSbIbr2pScoRwKyIYeaPVNVSeWw0dbitdHCRjL/CYqNjxc+nMBlJ/XZvpb2kHGam
zFyB9sh7GbmpWwlpDhvfLUTb0PckcayTEhQPYxa4EfBVdfqOdaqHBQ4KeGJiog7jkjcNPXBp4PFAtM7mq3J81e5n3DSNjQOk43druyfJS9O4YWjxaqk39rqDGQqHunr9
Kxzrje/F5wU1J9G1vZvdXwDgASXik00LHjocs0QsRMNAyaqwkAgzq4ApJkwTRqQM1VJ5bDR1uK10cJGMv8JiowpRjzp3eAqogEJZudqvO8/MXIH2yHsZualbCWkOG98t
RNvQ9yRxrJMSFA9jFrgR8NOOH6qI0YgOOX9t/ch7MaCSNw09cGng8UC0zuarcnzVpG8juvlWEtIQWqN3OYm8TbhhaPFqqTf2uoMZCoe6ev0rHOuN78XnBTUn0bW9m91f
nZ2bPqw1eUEzUTkkQnO1dEDJqrCQCDOrgCkmTBNGpAzVUnlsNHW4rXRwkYy/wmKj1ZMhar/1WZMK95yMOxpFo8xcgfbIexm5qVsJaQ4b3y1E29D3JHGskxIUD2MWuBHw
RWFmHgh68ExdJ1znzavicy8xkZyqNAXhCuc7grIB49JNrOe0POlmnvEHzG3DuAc+OChwhrvOT1+LtITHLffs5YiTzaeBQzdz2bF8pd5cNDLKiCbRJr2HgYyrX3ljAm2I
oFN7gHeT+ZseMhR+qjrtIoU2knnEs5OCk04qUddxYB/exP/PDYaK39CDcx/wIx10MM0UPyBALupT74JVMyKeLMqIJtEmvYeBjKtfeWMCbYj2iSZLDKheHdxeEn3nPbl3
1EUTgxCJ36b5TQOV2viBgu4KXaT+E4dahZ2DC7o0umDKdkmhOWd/n5cvNZX5BNjtXPOyDk3IC0mk6GbfpWB41DLhO2WUxhU4yxGZMmgUNXH36CaiRKboK5UYl3LJ7zx0
t3+eq9qpknE5Kp4VpkCCbFzzsg5NyAtJpOhm36VgeNQy4TtllMYVOMsRmTJoFDVxDNA7KqoFWMcXMYNA0WpFUpTWG0aB3BtHkEuTpQRdVQBc87IOTcgLSaToZt+lYHjU
MuE7ZZTGFTjLEZkyaBQ1cU3mzPdd4BsUy93gk+8I6WFsyoZ1oMsVikl4fPfhY0md8JoSnAHWaUwuSVzn5GP6JOr7r2n+y5s0zaFyglTdRxIc4I8bBRU4fq0V9K9Lk2hT
mqdMwR0MEKpM063cMUZhlcrUB/ytmPyswYjhbwjuAJqmesbmOL+i5BIjvtn3I+gpM45djlhp77QHgApCsFIShCFFaLQ1EVGN/JZT4UVOMydEX4DkrUNEzUikKvL5FwLm
3/l/8akIHpwx82+l8aNJvdMcdZjaLkSq2bXhn00eTq0XKd42S5UNTCdTd7l/0WXHveFNKiEGHU/LWvKYHs9K2dgxKvyaoYEwPzhNQOE/q+zsAF300tmjyI+L2k444QJ2
q3/imk8dTOTHmV3dj5tX5W7IfpunVZhrx6jgVU2gS6/MXIH2yHsZualbCWkOG98tP9qrET6eF7PH4vosV2V1J3LdBDcTKXZ8KfewW9c8k9Sn3CW80K28Dl+6xhv/7cZY
2DEq/JqhgTA/OE1A4T+r7OwAXfTS2aPIj4vaTjjhAnYkEp5zMfZT1hbf6NKcDexRMM06zAsD2tJ1Gn4dkASwNknMno60xbMMDpduPd2NkdSQL042ZKgHMWS2e796lxG2
gpZBSzNKBNXcraWGJROdJ62k4aLwcekbHiHWKN/pt2aFwAYU0KibJ9HvzaVNnMveFE+1rTBAP1xVI00uxjlcMz9SzSummDgzl3h21gExybUNZiIDoDIwToWdxG3qKjsX
qmYH9Uq7tL4DLSSHqhKTG/YFamVOfuMhc645F+SN5mcdxy3+MIUNj5NupjXeKR3WmozKuqkViTWKEFs0tWudcKKLpsBWu8O/ayZjdJtoSjUdG8ehsZXZRdtBw+vytX8q
hcAGFNComyfR782lTZzL3pLNj/VzF316t4Eix1dkct+QusrBEVuzjVdlwFWvfUNvoLLkqzo80iqutKG/oMm45ZFO/bv30Ym7s8s2vG+uaDVnxfqYIyOYnnbj3aWnRs6Z
6XO1/YppDLGicqU6296LO7zA6PXm2nPB0s9oYACUS7sNZiYDRIqEQjc9hKDVTBl9iAUR1LGetLbyDIPCtcWFLIw/9qE0bCxw363OXpvTHI0srBvwOnVXOa6JSwqdWbkz
3VmksQEKxYrogZjN1e3hrZW2gSTMD3+iImi/JcpwaUhi9zOn3PacG1bgxUmgbVBhwkByTZojkziKZXoORqK6aR+6rJ7Pt3a6Gzq/szqkCFvWdaNZJk3lMwxxT5blcT+8
CcXpb2GRrFO7e/wF0kXR4S+6NXPrsS9R1t5kboLMOhYjPlTJc+aE7PSzruqztFxmLC5dQz+p4/YgDcR2tmvKSAnF6W9hkaxTu3v8BdJF0eHEpMLlU3HvGi8vEgZaR8k+
aPz5N2F/CFsHLcHDNGxY/beTYF4wmhOT/pEnJGFyQ43QB4BrMk29YZeA8yBTDIUFZOXdcRjzbLYuU0iH7sGiIbmXZihz3TlxB/gRqbGBlqXymx8iWpuRfgfIuUB4bT5J
GZR2xub1d1sc9su6tWXPbRhXgvLe0SV4DMRXee2/Fx6lw+i+7TVoaBHiCNWvoeGihTONw6IJNb+15hXStSdG5GuYbSGxUB1H6tBvFTaJ1/YbzeIEn6dXgNiaApsv1Lbe
boe/Guo/QoJqgfu7V6OOffXf6ERKmWyjW5o4O+puJ2Yh8e9wrbiDv3A5RdYlXMRUm5Xnbx20WECZqicp51hpnkVP27pqi0WX5+i043ww9hgwLELNZbaSjnZh5Ked8J4w
SBOQesHmVZqBO4LfgOWcEhlIHESyk4Yner/E1nuE07kF8rwqS+stgKS07ZcCw1awymmHUfqg3+GFowhlaF84JKlrtBX5gx6k1p7lDBBK6vAfuqyez7d2uhs6v7M6pAhb
sS8cASzGj4ztvR2IaXud62HAl/Twbd71hyiHcjxWjPOnuyD6UaoUlCnm5K1en2VeB8Ix3PRfLXqJ72rtTRgQo7LNcim9ihnZ31LrTMUeXSGAfRXRyMwuoDgdKnwS5rS2
/k4N+xS1XQPEQXXj9ZPag7mvl7QQ+7b2aMhbItGElOolrhPCZ0++E9Jm4MHMHcCWiCezA71BHdOhSObaTIhU87ClJQaObMdQgBGrIL/wyOu2binpSv0rIEzzPDn2zWWh
h5DQ3XSbvAh0wCRiMivWWMEFJDxtCuNN5QydsMVvV3O5v3AQUZVLkUf0wk83vvLEQ0vekNgI13b+cHi6w8qIVfblgCXYlYp42JPBogKYIkp4e4vr1yuPGPhdti8Kxgnf
JtuF7KUASrRjbMZewYMKIw2VPTwGl8etwlQb9tcB8S6Cm7AS3fhnyv3vPbQZu6mmc/QBfy4s1n703UqmBVj1BnA7WFttYNVES55AMifDFNllE/IpTiBoeNKdLlRgtJgF
auNYhQoQL+nC+XAvO70KBgz9bKYVcmL+J/eUpOmKdziX2a5+4EzD963uZc5/3KlU6AlSfKXjk/ySoMCIBPTftCQD5OEqqp1D6TKlk1MEwpshO8uBTz+vy3zgIe0QNseP
JAPk4SqqnUPpMqWTUwTCm7+TKwJPvCcAm+PaJ7boF9kCOrAuHVn6t9v7Tzk2HCQrMpUjjQ60V2nXkY5MN247kdEyvqBV09Lgwmec71Yph75RHyZdY3sr1xhzv7vi0S6B
JsV3xmKDATfouyPvsAmfgp4IPVXg0OjhKh2dLCNGam17aNzBUm585CuDtg+hffA6AcTvF8gwooMKmKArv5m08DoehRXQM87rIlkPWZ9z+gvGzOQZZsXH4i3fYK+uLg+c
kikicTixje+niKPzA8hK3FgGGnrde3Q46YVENyLvX0DwCbUXa76PIAW1vrnZS91MYnD9NegiGooOXCkTmqo6s+BaeliaO+GoZF9REHtFssznx7hLcHt6FLJhxtObKePr
YdmcAqjnHV9+NgcZYS+qiy3Q9zckwBapNc9YrkLHiufJpynnhcjZFmq2AhJiFD5DH7XKnwS+eQv+30FXqg5yurqtTgABgf1h90jjSmYK8QbeC0AqoYVRhrzEZFCd7jZS
qjKOcI9gPfYCLPRjFKHvR2C2xmMQPCwc1Kr4OzCnOS6fqVFkwNibaXqp5aRl+ucTjjBQ75PEGCAZy4xAQPPuZ22S9yV2Tg0TPQve6ggf+B94UVgQc65mLsvpr+7e88bN
961Kjjok0iHYUyDIOR1Yrr18HfrY2CXtwN/0Ih39bGb8CvFL9nXrqXZvAioIb0/7S8dhLviyllgQw3kA2eKs+a+bnQ1Co666pKJnBPM/Du1ZxAO1toC4FAOBN49pt/qc
dJALm99oJlbWIUAK7CpzmK/UFbKCXPr/rxx/DATL/GDJ+crxX5Nkk9DoqT2fJmiDgIe5AJ3Na95E04g3cZN4TfaHgh6D2RfqPS5HUDIh8T9wjeZXcIFrutFp4NXX59Ey
4tfbohEqliyvQ/VLBvYnhbPqzge+g22Bp+dJaQJvBsDyvmZz4yN9O+15RfQ2gpzMXPOyDk3IC0mk6GbfpWB41EQW3586W/gOvmnfO58sVZ4tmY5kDygoEvwE+SriYkoc
GvrsxYmy1bezQ357ILAqDDFZJHm7e78hC0ZjLe4q6+5iq0ya44oBmX/GToOs6Y0ZAHTzE/M3DM4XIMIEr424t9wPz8YEGFoGCQsrXZ9ValFOGND1zCNp/M7TPcPCht/a
VYdnCuzy73AtTQiRVs41/NwzA5ZWs4PVUk7dJSuvz+yaIj3frYsws81ln2baUsNG8YjXWphvdKjibu+xVSDtpHW8eX38KFJxh4M8oTs+Sixh2ZwCqOcdX342BxlhL6qL
7zLyHoIwy1nSr/aexE5ps95aQt6urgtj0QXznq/S2z5cMjdTufMOnj2mRPwJV3k3oPejuWTbTvma9Hj0YVw56UNPo7VE7zEweS0fMj6bZ+P/EpVm2t5pDH+0KaXMLopd
AuSW9vKd9JBJplcCnjtbK0Lvxm2gwhpbKV50hz7nZJzk5c88MBBfmZSFp9dTUri58b0qqSjGDgcV77iDxmUsdK5mHxemdU7ceglzsywNVKXDYo7A7UfqN3WNTURpwaj3
bBAKYYZoMuVDposw4NVYQ38wBTNTNKYFHB3PgCEsnjX5zDESU9Qi15PClxfLXkX5DJc27TF1kHbbK+byo/nwaGJu4OJ43r/pgsYnaHd3zJJQtBujPI+t5rtAQzxvEYE2
XPOyDk3IC0mk6GbfpWB41EQW3586W/gOvmnfO58sVZ41iW4FzImSY1WiUIak6BAvGvrsxYmy1bezQ357ILAqDPlDPhr9AJ9c+QWadGZBMqdiq0ya44oBmX/GToOs6Y0Z
VEdLnnIIBWrOydAj13KuzcqIJtEmvYeBjKtfeWMCbYiwUMXej5HmBGke8IoEq07oZ9mU8SRMFQ9gIKnPJ+04OgiJhjuCuZzHuO0/ZmExXuSL7/tLHUPSEUkiHtDAVJd7
UlBYGNJSV6vyT7bPRhsdaONTRP4LziXVxrqrOgc92AhYBhp63Xt0OOmFRDci719AB4T+SKOyceAOXc7UJOVokpUvsBOX6tkCc789p8A0zlSYrVupKZv7UzB7rr6s+6Vs
AcTvF8gwooMKmKArv5m08MVb7avDHQuuoZq4xWYqm3L8CvFL9nXrqXZvAioIb0/7S8dhLviyllgQw3kA2eKs+dt/2NBiWcJJq0yUCocCX2Ni2oKEPiL45y88aYXW2Nvr
kWqwFva4erWXBR1Z2yEHCJRsEC3VGJytONxDNGbiyAckprrRgmofbDxvVQRsZSub3A/PxgQYWgYJCytdn1VqUU4Y0PXMI2n8ztM9w8KG39pBW25EF+LAxVsRKHfDAMbK
5BVlBYcwfiP9JljaIGcIQIvv+0sdQ9IRSSIe0MBUl3tSUFgY0lJXq/JPts9GGx1oq5WjMsBihkvRgD6cPFSPGlgGGnrde3Q46YVENyLvX0CAy9toAyXsf/3mhfOtLTXq
pBzUqNbl4Owgiq+8uIMlfV1ie+ddM69EGsQ2SbF8auH3rUqOOiTSIdhTIMg5HViu0wvEjE1wyQ86jPQmwS6gPNv2yrZbIQCHY3y8nboRbUY3iAK9zDdqWMnPX6bAlnlH
IHSOCXUcGXRw3NaWg/K6kBr67MWJstW3s0N+eyCwKgwgyB6lx4o6ZfsFwSPwVeCNYqtMmuOKAZl/xk6DrOmNGZVtLoz8JEbsI4RR6CS6TADKiCbRJr2HgYyrX3ljAm2I
sFDF3o+R5gRpHvCKBKtO6HnjVsCc4ppGRmDVV+AG0Oh/LgJsS3Lb8iYDEF4gHyK5/wCw8Z9KwwNpYlpQeXe/vy0I3sSM2Th/IybHqzqDBi5CYOuO03UdPGqW3oOn5jZK
b8918NcfoUYwWTmcsqbTcbblxf8UwL/TRURK0NB4tyJezh8DC+e2mJtBar7Yq1rl9AhpRkVDG1xSC2/f4LJ/B2Ju4OJ43r/pgsYnaHd3zJKUz0sUOTld6Z949CN2nQWI
W7dPjq/7jzHvleLIgISEWlgGGnrde3Q46YVENyLvX0BDQCMxLYPuejS3sj7ocBFferaMep6T5+iQeNZY9KMyu9DEj869zF5rMBOp/Y5qptPH/mlvhPoPndbzltRiMs1z
6blyApdsKqZbZoWwlJQtH3qyqcpUVsCINXgmVKejsUIC6rfHlK5fly0cmzdu4erl+Pi1AFoH/6bH31wbC7139dk0xTz68oe0P7D44LMBBO0mxXfGYoMBN+i7I++wCZ+C
GZR2xub1d1sc9su6tWXPbdUR7xDEra8OesYHPacT0Z2/yeF540gSCzOngDemuoXA612fT7RT+k/WQrAagB+5ybfXpze8KAJVqYFEtC7ilC+FQrVlxxHTrma1WIvDwtmb
s3g8u9kawj+8mpGWlANQ2+WZYe3KbzPKOZ+fBOGE74HGayNTfgw+V/mMnJIwqU4cKLdhgvm3UqAgl3WJoLDy89F6DC46HaVxNMmYzat8+fmEAMjww/k+ydsuVhDPBJ7T
vuSHSe2SLOg2E4BdZEw22lMArvqfdj1OM1u4OuwLpvrpfTg3We0ea27gMOoBM05pWAYaet17dDjphUQ3Iu9fQDBwuC0hcOz+rfwGjx8CCahBMTyuY7xkPU+8NrtnMzLJ
UTpy/FyqsFH2FO1cZkD3Snq2jHqek+fokHjWWPSjMru6AFzkarePup/6YDQtmbLU2/bKtlshAIdjfLyduhFtRsy21PlDVBvYXl7/ZxaaL+0UrDk77cfteA79vJSjhmZR
LNvVYRZbrBj6zSkoPGiAr5QyYJ9gk5rGiR9EKRi9iUFTAK76n3Y9TjNbuDrsC6b6lrHtCFE0wlEVqTrwnjwG7FgGGnrde3Q46YVENyLvX0CqPBTp34rdqNJ1Rgg9pKqm
WQ67rQOPunAFlArvM7HhKhRXKHN8MJpurM2b/17gahtFnibTU6QhBx+5S5wtNH6qu1O+I++aWNe03MS4ZDtEsuEVeYBtHot7eYFbO3lBiAFrb59C3lKcnIpeI0RPEpkX
p9phxuYz6t6+rYDsRtdDboQAyPDD+T7J2y5WEM8EntO+5IdJ7ZIs6DYTgF1kTDbaUwCu+p92PU4zW7g67Aum+mzngB6IZm+fyV5C8UgKFRtvz3Xw1x+hRjBZOZyyptNx
L00dClORFprQ6zFrqBxcZ/XUZwawDxiZp+BAodhCo1vwAewxC0LGRz/WZPIPK2/NYzTylLNIZrU1ICSo+xTWfcROWIPqqK6nnXL4mrsDCJN/QXQAldk/itQXYx4BVOdV
Xlgc2AeyiBZCKom810U05Jwax4jqIWDNw3F0+f95+XbJjGvFcST7EMn4DmkssqGswnEt9YTR+4YpvGlEyRquPmJu4OJ43r/pgsYnaHd3zJLx+y+TtomDkkUUhVKxOaSw
tG2m3FYQ9JxYqHVEDSHPpKE/BDWGc47iBePYe0/9mVYB6lOdFRqfT2TIA4o3J4xE1UmthPARkaz7pezGesV+3n09ZnqVXtM9HTvgiAICZ7CMJogCCP/b4xI/jvKx6iDB
qyClerOV2KTffH46H+fa0mHZnAKo5x1ffjYHGWEvqoug4m8MpvMTrp+agV1WlxhY20zzQqpU+uUEifcwvtf/sP2YIHkDYy/RCCTjZnpsuK6dG77qT0pL/25BPXQ9DqBy
h2lTBLcoRewirAaNNr7NFPwK8Uv2deupdm8CKghvT/vlPpnYBcj92m7Yzs6EjX2DSO+27igbVuqqAQ65L9uaOLmCrj2RE+0hbJllu18Pxtt4VWMvY9+wbp7oLkpgtP08
4Fp6WJo74ahkX1EQe0WyzGvUtq5wcvhxLm39TV7ddcDbvgMINEPwcf7e/tubne8PYOKSSGOOl8FSoUpX0xsRLauUd4EpaP5iQWlocZPaMsld+hmW+andBn7dF3juH52F
euYsyRojEq/8DF2CyR/+SQrBg22L7Aqu2KI6TLwxRtPhFXmAbR6Le3mBWzt5QYgBa2+fQt5SnJyKXiNETxKZF0HGiZrL4m2OeYF7wb1z6fWEAMjww/k+ydsuVhDPBJ7T
DfZUysjJ1NyiHx+VmeVhSfetSo46JNIh2FMgyDkdWK5fo8eH1mJicKpcjs5nv40oJsV3xmKDATfouyPvsAmfgvzmyQ5CrjLjGMDjYYshQJz19odiTrVsBvAAMS/sjffX
4EbrQ1azvA3FJSGuw+C46vqU8hkCQNI34Myh03N9mzbFSd2Los5ywaAGfzOSde8fqClh2gBZfYcOROx/RoLPGUQW3586W/gOvmnfO58sVZ4DpXhvGD0LwYls2xfBGqSn
yvhVAGHHiE+eq7WHFRJY6wAihdYX1SzpZBDyLN0CpE2kLZYL6uR6f2MDl/DROfp5Qc9QrsKOaijhLuQgL9s3sNv2yrZbIQCHY3y8nboRbUbMttT5Q1Qb2F5e/2cWmi/t
sBIBqqmEQqJUhsrdvsXLvIQAyPDD+T7J2y5WEM8EntM0J8F82IjDCeLgpWcQ1ztg961Kjjok0iHYUyDIOR1YrqoKa/cUnqL9uyhHIZMiNjUmxXfGYoMBN+i7I++wCZ+C
/ObJDkKuMuMYwONhiyFAnLnl/NB/o4G2xEgdUvNSC/wHQ10K/sWHUz49dZX1enIZ4ciKDpacDFtN9fw8G3qfcDDDqAmfjK1k2sDcBT9bnQfLKmbzbwxkc1CtF/lkhwhQ
UvGZT0PoG8FqPaEC9eivn3+h1AubXFHSNdxRHAWmxsUSa/eThv11imJ8yCU8icruehxJh26eG0iu/A7AE000wMVzDO5KtKd+ibwrn5U6xlWmQS1Me/LOuEnQAqI6FYXv
W8fMhQq4ZCXWmBd7OMO2eisc643vxecFNSfRtb2b3V+Qcw/mYsBjWSIUAIuFFGiq/ArxS/Z166l2bwIqCG9P+x2cg79mx3l+S4DSmudXL4PUf6KMCAtteyT8ci26Xplj
eraMep6T5+iQeNZY9KMyuyDpVcwJqBBfqlS9TuEl7NRozOIjrrGS5B2OX/mDcX9531UP3h+S+PJOrlKjdX7z2+oRF8IH9xTSSMBAlFNs4KdFha3BqO/K6nU5OevzxoBQ
9d/oREqZbKNbmjg76m4nZmxP3DIUPzZR/cap5+Ns+mykLZYL6uR6f2MDl/DROfp5+tXHwpyNNCOAxnMHvABqYGNE3Q7FT2pd7hcimsiiGf7HfWojvrM/wXvjC8LipbjA
Q3khgLg497t91cWmpYIiVbRtptxWEPScWKh1RA0hz6QqEgimWUdLnWGKYVZPSE4INNzXYOabUIydeiSiCh0wRp0bvupPSkv/bkE9dD0OoHJl2mt5153CYUqezAkOOPsF
zhhICemm4c++A+eKp+MMaiVBLY80EXe8En26Fhz/wdht3o6YKyn5MUJ+MNPiaw7GJsV3xmKDATfouyPvsAmfghmUdsbm9XdbHPbLurVlz23Ms4/W7ABi3jXc951Xl2zX
s+rOB76DbYGn50lpAm8GwJH3TnQvLDzIMltOROcGrQGJo1uMWgoVBZoQI95J3oxm31UP3h+S+PJOrlKjdX7z2wnJs6AIDWX67qYRfYLEzTUaN8VUf1vcyWeYxahthnWt
6QOdOeia+AF0eWdC1ACaUNuZJndI4bQI6M9sd3ShGMpG0ApRjLCd4PgaFzEbTNXupEnbFB+ubSMQP9sUGZbjRt/TIyWPg03JznnB/AkGQ1u33P4wPGqba0lozzMDg1jT
j1AnSXLTNSF9DEw7RUMeig9M0diUUth7Umdt0QY6a9PfVQ/eH5L48k6uUqN1fvPbeuw81V6Ie92qqIhQs2/stR3mgYkv0pCDymmWXQ+EwdvUgcyDVvDwzjtIkqkGkLWp
qxtknDJtUqX9hYiLLWUcoTfgQ4OxB6r26o/8ZZqS6LV0m4EEG9mVJ17dWE5OAOZ/k7WHqsUyLMn74LbAxSEa4qd+Z47+dSokrBU1fSZE1x5rjkBAT4K9Fu0Qt/XM+emi
eFLEFgxhMNgk9gTBLvhWQOu9iSp6hfStMsJxhHyV3tXhJ/GtpzphEEFLy7/0nBZ9qZKlq3+DX9dKlMfzulBc8agPeRSiiiBSLrNM6L/oJvajEenPzO3tjOs0cehlNUIP
qVu6MnaBCMysuW8+bF32tCBp8yEWG4dufaL5F6K7WawFjTfBTsqe9BM1tHQPYURk1cgtwNMgvuQRs/yhfkjB8BwGM91Je7ndQoJOhBSVO+cjNxyGXxDrgNl28BoCebbM
x7/4b2NCIuZEKeOqcNz3o5zY9XYuQOKfVQvmPDwrecQ3U1Vptlhb24CpO+NUK7/AHHFmLwr4eHi8nGNaFJfXE1UociUv/V9K2/+e/T56MiHB51hOD63lnzcz5x7X2MCu
J3yadE7pOT2Y9l9asRPn4FgF9GkqvI3T532KH4N1qB2vRCaMKfb8q26yR6NXzAUfLxJt+lUud/jHHJy8uOPU/6gPeRSiiiBSLrNM6L/oJvaI6dYtGc6N6xGFXGW7F/DQ
1NmhPqDRLNcGg+OzsAiVPhRiwHZJEJ1ypqqKgExMB/bp4hHPvXL6044wcAOCMKOWb2c/FhwgFm76cayrLhJAP2zSDM9tbunqQe32suFmdCyTTd9zo9gXac2imlfVhkL9
fIc+LFYiABY4ZQF5z855mLGCFakWnP4Vz/w+Gh9cyi5z85KGOCdgMGccuMhJHaqR/YAgPyM4+p4KL4VJHaugyx2W+TcdZwhezt/d89Ty/mnG6sb6W+ulySnSp/E0BIwt
ZKEsrDLsaAy65eYaiu3MBjgFy7p2AZ9iO7hMJgaPzEBKLSoun8vN8YVEJXMFqGmCVHPvznLvsa87860LinhlSYsnZXY+8KIQYQ74qqtSm1DSU1e4W63JqbXbjhHggEba
b2c/FhwgFm76cayrLhJAP/dzimPm3b/7UmfJN0OyIhjq30qXqWFe6ZIjKsYiJu4FnmFo83c8IazQxWNbcd6dvMqC3dT1hgkdIOGph9AtLfNQ4UnBkDIrATBm7se0jqV8
+T2w9EQ2sWbu/l5M4S56BJGeUU4iECllVU2YvarbztYM7gE7AGYFG4Yb8pAFf2Dm/vvn9dbmteL/M1x3aiQ3YVDhScGQMisBMGbux7SOpXzQ5lfpdZziNvOhVjrj3Ma3
Mm6MhkT2xsI7GFqisSHP7v9+Iwi/SPt6VedfFOTCa2K8iLysP6xbnrIrKGJ7SCPd2BgpzMpqo3IiCSMNPNRaLxRiwHZJEJ1ypqqKgExMB/Z0pCFUG1R/Du0PKQwKFdgr
OAXLunYBn2I7uEwmBo/MQLZnoEoDU9Ejk0IfmQ9WrBY+TFICXsmb/VYbXBkpTK6cOe6kapocTXX5y0vkjXsQcpmueiAVo+DqPWi1+3g+vuPEmBPSk0KCZ5KTVBLjAZeB
PJzWF8qlT2ahBX+F7yHVs0ANyBrfaQOfCYSlPvxxmk8M7gE7AGYFG4Yb8pAFf2Dmi80oYW7AyAppAjnnNtL6yBCJLOS+HkbD+vejgUAUYcF+FLqUoYWgfB7tzHlVe3fx
8j1PtH7t74iLQqJFN4bVQDs+FcowHIPWZY/nMBcBQ17lsMsVULjzg1VT4Bk229jMlmTBv/Jsyh2wrXC7dMiOos3OqvbosFkAM/spQ1QrRbLa1R5F6uYLgUt0AH/9Dq/9
GYKHFdS0GuQhYkLUEvNgx9xW79ggHmK576Sk4cfLrXEH39EmOMVMnxKb/oAbdJxx62sdUJBGmnwIAri7z3dXY8uSubm2FbAP1BsGY+lvtQO8eMDU3kwq8F6AsCz++QZz
5xvZvaXfIzWm0lUDJAFNH5I2ShFO+KpOjmHATRCKzVGQl7R1G73J1Kx0A556GbKO6cVg6/S8FksDy0N+zK0AJjs+FcowHIPWZY/nMBcBQ16/W52X2SMUNi51jDNuSv8b
dJuBBBvZlSde3VhOTgDmf03ficgDsM3KiLrTnZZdw4I+I0zWPlMHWSZMRWYRZ204HmcEzAtP6wSVwuUCrOrzcFPwOFf40lQ2LzLJqN8XWhQDB0hKzR5X2Xg4qqFzz6U6
J9lyxuvwBLQhdy6MxQNGJ+Fyz+JlfL5iIkGXOkvCQRmLJ2V2PvCiEGEO+KqrUptQc43FJF+BWbFocmwhvA0w5CTgMk4XjNz7CIfPz+6cVSHKiCbRJr2HgYyrX3ljAm2I
5hv+l6hU29B9lbevukpQxk1LYgM9AnSljnX/4EzcvU2Lyr6lAMTJ9WMf+Bi1PTyVVqVXrcGgaMOJfWNHzCMZ6+lztf2KaQyxonKlOtveizup/dtG1HjVhLN+xGE047d3
Jz1MjxVV/HCqTvskm/mtyGePFjGOfzbu/bLM8i364ZqClkFLM0oE1dytpYYlE50n99pWHgy8TI7u5vLZ9799vyBp8yEWG4dufaL5F6K7WawgmkqmfVChLUn3aGQEZP6l
rNYQEMWcbSiwWe7mDu7LWEg75Ye0HKEzWEmbB55VD3YWAOWCELPqYw3s9eqzjt7lSnFYigBMVulUQAL9JYT7SwOo1sr8/HpHKasIVByYQH5JYySJWlq+qXWZJR8Pwqb0
ZGx7PaewS5jsXOzwENMZvBto1TruR4eZ1tECV23cD25/8FbGTmyEko9NwfApVa0/RMe0g7shdEuSAHNcBohXCeYb/peoVNvQfZW3r7pKUMaii6bAVrvDv2smY3SbaEo1
hXNXuCwdvPLv3euh+7IrEdILvtLImYKbqdQNjKCXwWVzjcUkX4FZsWhybCG8DTDkoXXvS3wxDP4SYbI++QUVxqkEofYL2Vt8CT+Zq2w7U0Tp970xIkM8CExTRqTEeRQ5
SnFYigBMVulUQAL9JYT7S8JAck2aI5M4imV6Dkaiumm0ouNgomzjPv4xDxjaN1sjHAYz3Ul7ud1Cgk6EFJU75287Zke/GxiZJK1MfihgcY8gDvtYVzG7xwtKpSL+MNii
lkfiVouvsklfgOyR/fbyHmePFjGOfzbu/bLM8i364ZqClkFLM0oE1dytpYYlE50n6yP2dMWIBR/wvUiUeh/7fYsnZXY+8KIQYQ74qqtSm1BzjcUkX4FZsWhybCG8DTDk
emJo7//OxIByLo+VTlkjE1bjsPeUkDv9UO3yj2H0C5yixe8ZJPYoFH9o2EI8M5ENehxJh26eG0iu/A7AE000wGye/qnUSClHmoVadCQJ1xccWdHPYxB18uMkj1Emgh2F
u88f74Q0xapWqUSTryYEMkTb0PckcayTEhQPYxa4EfC9j4b+2WyrQpbTopmuMgK6V0qtsc0oR7X06bTRgur/mV32DmI9Mck5+/ph3Wtvdj7XtBIuo29rZQI30HT9ns0l
q3J1SjMH1k4FLkVcmJSM3RwGM91Je7ndQoJOhBSVO+crHOuN78XnBTUn0bW9m91f8NLwqB3K2vL5MzA3pzbolJZH4laLr7JJX4Dskf328h5njxYxjn827v2yzPIt+uGa
RtAKUYywneD4GhcxG0zV7nluzcM9End/yld54NU2qSijQ0tcWUt86HTM50PupoMYc43FJF+BWbFocmwhvA0w5PjOggMTnTOANd3zkh4wa0dqhLmMpKk7K4MJpnjub3A4
EiR2gDb0d/y4CjT7PTh/in45kPdRv4f8skOKw+Y7HRkT0owtUUO3drlx4zryJdPwtKLjYKJs4z7+MQ8Y2jdbIxwGM91Je7ndQoJOhBSVO+crHOuN78XnBTUn0bW9m91f
J8y8tdD5L0ftGU4gBcFTwkLZJnxFLR+05+2wLmZ9l/tECjsXJb1HkW6rtLAsWEGdJUEtjzQRd7wSfboWHP/B2G0pdElQ+CA/eQEVJb8uZk3Hv/hvY0Ii5kQp46pw3Pej
u88f74Q0xapWqUSTryYEMkTb0PckcayTEhQPYxa4EfCaJ0m40H72SbaB7mc501qHWAYaet17dDjphUQ3Iu9fQA5MhQDRvFuaGZWQgnm8BLxVCfsglt/Uc4QUSxecuTuR
rZY+XdSkH4lY6omSSWNTV9NEKVMacbim6wAuo0FkOkvyCnzYr6/pXQClC2C2PNIHeVvA2+3eVAbws3VQmjKDuiO5c24CEo9fOl0TtLIhRI6GRTy8fKkaJ3S+Wm7WTxzC
dysZgBq/QaFXLj5PB4EQwQolaWFRjC3BJ8GRnajb5fzmjYZGTPpx5fHkDH12aeTGjXW1QcpnKZtQ3fqY30dVp5vcR1dZbqYcU/1sbWGAsF8xm+oZsSbUW+jr2g7j+WMi
lkfiVouvsklfgOyR/fbyHrhKly2+93psrLOhbt2R96dT9lzAVlJp4jL9ic6fWHtrNplpTDK4lIBf6rIUe9FOVSc9TI8VVfxwqk77JJv5rci4Spctvvd6bKyzoW7dkfen
U/ZcwFZSaeIy/YnOn1h7a8hCHPCheslXMUMukcrCvmcbrxcGe7he+qeufjGLZjeIeKFt9AgoUGZlAKIsRIF2Qw9j7PCZPvgatTifBjuV941PXeymvg9/bL7wb9A6EDAm
YAl5qRUKcux0ZzUQsvMXPlFHc8xtHUVYH5az6Bo1wQhCbx3DvkQzB6gGOEg1jtBYrZY+XdSkH4lY6omSSWNTV2dWjGi78idoW9uXhbVLjT/MB+9cadiOnkTQ0lTocvF6
hGGPl6Cq2k5SfVx8BCf5Avyn1KOhysesLtv5hC9TjqS6Qh0IRWUf+aWXV8DdowRy/pENDS1ZbFXwzFrnj/h07OaNhkZM+nHl8eQMfXZp5MbmUIzTZIC81+GPhmeJvoh9
BSS/vktns5jVOZzmpTrvVYTeC0hgYM2ANwGqrx42AyOrq9RmpYrYbtZS3UzuUjoHzEUIMAj05X0YRI7ZQ2Apl2OhTaE8BmnCtezcEt23D03qQyRncurkRGnYc/E/NvGs
kaX69Enp7Cx8xhBMiqW9NqStiTsMr4V06D3UL5pFaa0ysJ25GTPKWsu5Kgw5yOCnb2eeGVJ3ceTQ3DoyHOo/Wit4yzJRwMwbtPp+vPYF5BE0bgRG10JwQzuu46ahyNf0
KEo2dWGEJ6HycYwN6I80dw3LpqN3sex8+oZ44gR9q9Dqbjh6O/sSig7jjS3frL3t0nJzBMNJ1R/rn5OCXu9NLKoFvfpKw0kziEsXWgLK4XFsEAphhmgy5UOmizDg1VhD
GFYfdLtjZMDXlwWUIKHiveP9uRzUEnHTeJuWizEiQUzbvgMINEPwcf7e/tubne8PJkYQCLjgKnxTlersH3NsC7Si42CibOM+/jEPGNo3WyP6ADLJbFdBaUdz4Cjoq6XO
cSSLsEFU9EQIkYGT2zoXu4jpFgEfttsXL919vwAY910juXNuAhKPXzpdE7SyIUSOFokiG0igr83E8kenI3eFyeMEwOTFvGmAFhRj/ayuRnsdDnDV4VvQlhOsqttR41jm
n03a+ss7C146NmK/FakidjISJkZ/79gDZFmBNtk9qGi0ouNgomzjPv4xDxjaN1sj+gAyyWxXQWlHc+Ao6KulznEki7BBVPRECJGBk9s6F7vB0FMP+zosykyCC0XWLW24
YAl5qRUKcux0ZzUQsvMXPqzjZgR/Y7H//czrtmdid5FsEAphhmgy5UOmizDg1VhDJM3oJIu5gmy9p9izJCaziOaNhkZM+nHl8eQMfXZp5MZ6jO3qA7AOv08U4QVlxrCt
p69i7qjPkiM7wd8xO8b+3tsmY0BHd+m/6eufJjOlO1YNl8gNLPbM8AyjBiKynO1tI7lzbgISj186XRO0siFEjhmUdsbm9XdbHPbLurVlz20Qpc5Em1zY3cHbmt/pt8u1
e3yrtFw+gdllgfzOQcHFevFsm1xRQs+4Kt/kJpxmiTYC+FO+WzTfdDz3nS/zmT3uKmoblzZF9fi8giqcSOhB9VpXvilHq8/3or+u8OyEF3Aivd2N3DaA++kSca0KJLwD
etfygzRS4Wv5rAmruCljjWwzMHjRc61zJJm2SW/vv7JWPDhpe4Kexq8Qnxt+fRpj1fLc1Zj3cvHefv+H29SubHuTccXltOSzw5ShITFHqKrrKatqohmjJPWMzMTVF3lc
4KW5iWOpPFbfxIdsQX6RdlpoI5LHvtBep91ofqGfb6wr93VEsbBMkqdGW5pAhW31cgYyKnXcGPnun5d6d0mNe80UmJxS//aXL+6B5uIEP2zojQpj/T7hOm/1PaUHjPwH
L23lWB/TrP+q9Ztl/TXjZj/amu4fhMj7WPFqF8vHAYfaEwpntNvPt1yqyJOCvmGv58idQD1lZt14QvFBSamfEk28PlUiNHIKts41V/JjjXElQS2PNBF3vBJ9uhYc/8HY
iu7wl20zJ+LKoGd9RK3UxW7ncLBiTTGtVlzMi1r4pUWmZt8XW0UBNA3PikAT6QDyzE8gM3ZxYLlNVA1bEgCiz6AGc551tYbuYlsnRRbLcrQgsg4PXLogdu9DP+x+2EbU
ZdeUuzkLBjeXRCsJYLpduv30V66wF6qdNd43hTszrxyQ0PSc3WkjpV0VOA/mSK6CiS2cGpy3CllLY1vllopdcvaYsIGffv5N8A8q40a1fNSgED2AkrtRo+DC2Vuj7JuP
iKnFoURnRvLoSl8JH/TGhCGffKrKJPF6GBiUoVEM9NDazI+RAOr9d5AmokykP7PMWaFzyF99kpePBbWVPNrbEneeYPZp+fdYyu9EkfFHbIlu0NbUfvhlpW/s6StCJC6W
EiRmyFlI7fWVrvsEk7Z1FgGj1P7m+HGPKg4cS8q5gqZuTn+aVgREFQoWqdUOvLdv3fdyYNKT1Io2V6H63wgKobhRfnuk1a7KAvNsm2apf/BB98ZwR7PgJ7voYCWd7gtX
yogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUZ1AB+02V5BXdjMlgfKRVsHMuHGaFiqC0Va40HOdhiySzLSwrQyZi1/cWS6EqLaN338bUaFrrUWrJ3C8NEGi0zH
2IxgPx4X0/eBdEw8eySRiEDJqrCQCDOrgCkmTBNGpAyuLUiaGSbRvMiO2Y5sCASNAiINzVxRhiIGSrTN6PWs1u/+//3zFuBc6hpPyFOP3hyWYnCpLHNzGAC4XS62ftEe
9eAhsbYpcvuVPp86ImPIqn19gEBZcosw71mff8zTfJfpOQwmyrJONThm8bNO2Fti6LHUMREqEBXOZLt6guyLE5bwzClTy4XZndapCNNU+PPeBEehDRu5tBQw9W4ARUw6
3A/HQUAYHGYwc9euKnMf/O+Th44/BTRBMoPlJd1MJT/FgieKj3bLeSCOFOyV8tz5t0w3BgnPdKpADgobuDZ+ocqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFz
nJ/ke6EXREq9YL0GI/SkXGwRJGuzlB+/3aTi2zR/MO3Rv5n4W+QwCGZG/hQ4CIPeVMaUMndBwF+kwMksXvheRp5DxCzEkASNymFUZ4DxMUYTiY/nIHLUaG7nhQ7jQlgh
sjuddenln8ac5VYKnkY8n52gd7sS9grQRN9+GjLa5hxXavGLJ6DWVSg7vYWTRSGBT0AdSo0+Ioxd3pOapgecMXmXi0cBBNzIp1U7i75hqCC+nMFcJRniBj9+MV4li88z
cguOlyTEP3LaPcSElVlWBGi4oLzESENfX3xtj2wUKEDKiCbRJr2HgYyrX3ljAm2IdEMpVk0/iVLB/Xc8gKO+AyQJUjdB8uRmWExm8WrFdwHUsLylijY3gkKh/X990ZjI
WiozZBD53nvxqcPiINtO7cqIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0i70HRoP7GfTHaJ0xeliBg2Wy3NTGmkLbbDnI2+3pIrbdcKILqpViMAh92kTQwZ529
MKS9qjr8DhbiP98e3EH+StMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o3ea9yDxSSJF3wt1QQcMeY/UOzgVhr2GoovWyiZv7yByJscESQBuj93nozknI0ZC5
yogm0Sa9h4GMq195YwJtiFTpyjrT/nGj47Eokd8Uqh1E7oBqgUkTyQDTN8Kl7aOO8EdSPUz4/+iCZhpsB7CeFyHJYLdXEYCcJEEEwPiQI+NuPcqjj4KMfzKD264bGZmd
gRrInBgZD19HN9j5BZzno87kdbcVAiUyz7ljCbFNI5CflEwYHZwQwKKuv2jqpVYO5hv+l6hU29B9lbevukpQxlNsBzzkmI8VT8mzzaEM84/eBEehDRu5tBQw9W4ARUw6
K09CAaC+GdPoTocIAxv5eBzy/vYxc5wDFeFO2pzsq1pnE9PRDtnwCVnPJi7Ue/W6VOF9g7sh94P6znjjyr4gqsqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFG
qJI7YEbeIAYkNBFAqjXCBKH7e6XgzvuduYi+LZn7u0KyqEJyu3i4gKdJTpzWu/aCTNaw+g53QpRJfxKWC0Pwy+cDINPdkN0IRxIRWcP/qasSRqiVp9bf6hq6IpjBQBhW
Sly4z0Sxtnw0VPtn4NIa2mCAoeqsGCXzyB72PGVSnGp+OZD3Ub+H/LJDisPmOx0ZkQvSanyvBAlBVbKh6MPoQut48B4+Bk09Fg9hYF35DqKokjtgRt4gBiQ0EUCqNcIE
ay7DS6XVXYcYFc2rT2jws7KoQnK7eLiAp0lOnNa79oJM1rD6DndClEl/EpYLQ/DLIM/AlvMnyp7b1++Eh9RfUxJGqJWn1t/qGroimMFAGFahde9LfDEM/hJhsj75BRXG
sbuM5xjuyd3myH3AOqOAiX45kPdRv4f8skOKw+Y7HRmf8wPvZVcs+0N3jEMPJq02vIUBs7AlkTdVO5sdbY17dqiSO2BG3iAGJDQRQKo1wgR/lodsBscqqdPAbQkXGQyo
sqhCcrt4uICnSU6c1rv2gkzWsPoOd0KUSX8SlgtD8MvQZueJC7GqmVyxhdkNqLPcEkaolafW3+oauiKYwUAYVpzJPIvrIemSLOsF+r17NbpUoCwFEL7owHPR9y+0MRct
fjmQ91G/h/yyQ4rD5jsdGaB1uDZqewDNWmSw1fc/jo8i0ZW9YE28/xo0lLYLkHpYqJI7YEbeIAYkNBFAqjXCBBF1bUcFb7IWO/p955pUqLGyqEJyu3i4gKdJTpzWu/aC
TNaw+g53QpRJfxKWC0Pwywng564rQ9UHYyCLSeSZBhESRqiVp9bf6hq6IpjBQBhW4g3GhXDWW6dgddRYU5141AiqVzqYDVqOCASAYMPHNt1+OZD3Ub+H/LJDisPmOx0Z
71dCMIWBe1z6ZQYcPSesmhpfTP+ipNTNECc+nUgZh1+okjtgRt4gBiQ0EUCqNcIEwCPxXrQRguqcT1WD1pk7gbKoQnK7eLiAp0lOnNa79oJM1rD6DndClEl/EpYLQ/DL
LEG9tkZz7ih0UOnVipii7xJGqJWn1t/qGroimMFAGFbxgo6S2FjIiZAxtGi+DwOZgiErpBjMSd8XR6j8KvZWDX45kPdRv4f8skOKw+Y7HRnEpMLlU3HvGi8vEgZaR8k+
zaH4aZqWliI6V5x73u2dS8LAA8SMJD4sHLNJVt6Ew7+LYGtvY/Vs1h2pytLRB97EsqhCcrt4uICnSU6c1rv2gq2Jsefd6Qwy3BTLGnHfQcpNf3RUCPmzaE3QNwrVymL0
EkaolafW3+oauiKYwUAYVtxvP2XNaKMs6Ppux8JBg7d8i2uKIOe7JHQpwMhpIo7RzlCzuXDiTtCVhudFi/9xiNiMYD8eF9P3gXRMPHskkYjTIZGc9kTWzrYMDyDvnYgc
uc/k+OXiweAW5ELnA4Vm4MljTIfYsCq6sEaHJiunc2copYIO1NLAv81sj1hVgi//Kxzrje/F5wU1J9G1vZvdX1TsZmG/xjlD8L/OUTqK0i2JC7IMZSw1YTfxa19ZyEOu
1VJ5bDR1uK10cJGMv8Jio5Fe3SGfe+t89Oc4F/fdbLS7zx/vhDTFqlapRJOvJgQyRNvQ9yRxrJMSFA9jFrgR8D/+yQWpzwVNklE3mIVLoFOSNw09cGng8UC0zuarcnzV
EsSzcNPaHZ3v3QbrniXWrwbGTKeT40jgK2mkNftz9KMrHOuN78XnBTUn0bW9m91fFNhrSGCVVpYL3ESqjM55yJcxlX9YO+c3TxxC0LDHZG7VUnlsNHW4rXRwkYy/wmKj
89CR5KVNEaw9KqOqIkmdMLvPH++ENMWqVqlEk68mBDJE29D3JHGskxIUD2MWuBHwatsRNq43z+TIsPBtCPExRZI3DT1waeDxQLTO5qtyfNVKtdon1fV06N8NgVamJdxf
KKWCDtTSwL/NbI9YVYIv/ysc643vxecFNSfRtb2b3V8XRKkxIPoqpes/yrAnvj6ApSbIbr2pScoRwKyIYeaPVNVSeWw0dbitdHCRjL/CYqNjxc+nMBlJ/XZvpb2kHGam
u88f74Q0xapWqUSTryYEMkTb0PckcayTEhQPYxa4EfBVdfqOdaqHBQ4KeGJiog7jkjcNPXBp4PFAtM7mq3J81e5n3DSNjQOk43druyfJS9MopYIO1NLAv81sj1hVgi//
Kxzrje/F5wU1J9G1vZvdXwDgASXik00LHjocs0QsRMNAyaqwkAgzq4ApJkwTRqQM1VJ5bDR1uK10cJGMv8JiowpRjzp3eAqogEJZudqvO8+7zx/vhDTFqlapRJOvJgQy
RNvQ9yRxrJMSFA9jFrgR8NOOH6qI0YgOOX9t/ch7MaCSNw09cGng8UC0zuarcnzVpG8juvlWEtIQWqN3OYm8TSilgg7U0sC/zWyPWFWCL/8rHOuN78XnBTUn0bW9m91f
nZ2bPqw1eUEzUTkkQnO1dEDJqrCQCDOrgCkmTBNGpAzVUnlsNHW4rXRwkYy/wmKj1ZMhar/1WZMK95yMOxpFo7vPH++ENMWqVqlEk68mBDJE29D3JHGskxIUD2MWuBHw
RWFmHgh68ExdJ1znzavicy8xkZyqNAXhCuc7grIB49JNrOe0POlmnvEHzG3DuAc+OChwhrvOT1+LtITHLffs5YiTzaeBQzdz2bF8pd5cNDLKiCbRJr2HgYyrX3ljAm2I
oFN7gHeT+ZseMhR+qjrtIoU2knnEs5OCk04qUddxYB/exP/PDYaK39CDcx/wIx10MM0UPyBALupT74JVMyKeLMqIJtEmvYeBjKtfeWMCbYihwMxE2AHVTnC2UOYczdFt
d7kFW5P3dLTvQMORn7vyO23TFa5wW5gsAzJOgnxYU6LaN9TrbEqDpHsDjXIImnPG7lKbh9EN7lwc97Ho35jwjoYrbMx566uobBEB4EokLKoG/l2Lv0ueRUv92uDxdR6g
yogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKrNIuz5P/6n+zU0W4Q3q6kxsVKQRByGDQIIrBrQWW+c6p0x5fy9M8ITcNFAFVgTkIfzCE/ypZqavJ8qrUtEweu3
XIA6IN7aK96lFqPI7XaeZomvX5jRYBoyP+S0/fQvdRrASxl9VEBhpUgbNC/zmIYJHEtWIvD83khq2Yt6ymSRX2Ca0Ljd5eGriyCjL9D/ZC70CI663q+vi+PLu+pISS6a
Rdy5PvRglrwdSL+aTHC2TXfhVAV2dy9zisaodInfmAwV51tXjLbcMSf/AW0uGzI4HvCdZq+czYAXg8Ol5reAYkHc4QIkqPRIwrTppXiD6xsZBYUopuLNpWFxbc4yrTAl
T0AdSo0+Ioxd3pOapgecMX02msHhyGAcyZvVTmw5CwdLFVT2T+LoscguD6pNok9HhitszHnrq6hsEQHgSiQsqnEki7BBVPRECJGBk9s6F7vAgkmPjGDrWZ9z3bg+iKrS
9eAhsbYpcvuVPp86ImPIqnj2RU3C9WEk8zIsVxm9ceDpOQwmyrJONThm8bNO2FtinTHl/L0zwhNw0UAVWBOQh+dDIAyJu7m3FAP1jGhbX7wyzpinzexsSKNI9UWW2xEw
KbAWmvuvd8ilV1icDV9dy01Fq2X8PDypy9e1pLnHcsNn4QoHm3luxmY7MH2O7IMmYJrQuN3l4auLIKMv0P9kLgyXKoZBGRWR/PyJ9YAJCoZNf3RUCPmzaE3QNwrVymL0
xrWiYC43u26AAWvP4zXni9VIFMUCIbodJWI7MYsd30IHvi9svv2sIBtIX3uxjDSAyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhPQB1KjT4ijF3ek5qmB5wx
qUjMTPS9J1uVjYrA0qnoz5hWPQ7X/yoeIwRnXmEeH6WGK2zMeeurqGwRAeBKJCyqeZ+KFLwtGfDMmYbrekVCbysVimgSra5In2fQUEypWXBOMIr6t8q7SyEHxV39VfOk
WKxYHKySPn+8NepkuZ2mfwfjHCwMmsmIwx3KK9blikOdMeX8vTPCE3DRQBVYE5CHYaeA8HVsD0RSj1WQvO07IgEOEBoqqkgfO3BgnPoSl8k4rynSNkKO910BP0ILPGQH
EoyMTiT+Spx5h33PO1+Yy5SvK70Uc3nDR+4nGVTVE6BgmtC43eXhq4sgoy/Q/2QuwIgZwLJjzLxFZV9k7f1gr9Bm54kLsaqZXLGF2Q2os9zGtaJgLje7boABa8/jNeeL
zK/S5LhiBvAHc4X/K3S5iXyLa4og57skdCnAyGkijtEOTIUA0bxbmhmVkIJ5vAS8FRe8MsfaJ/3lhUEcM6pUCc9QzJxZT3F9wJOayCVO+QSa0pY/DuluUIHvmvQa47tU
OP8FoDq0i1xV19PKzLcyqWz8ECDuNb+dWCJTy1WrWqrKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKqpuW/zGTY+jlEvs5VC41/r
RGaQh+QnKXYFHTDKJU/xNZ0x5fy9M8ITcNFAFVgTkIffwc0NqB3BkuQfRGBsoTGBIp2+UGVxdzy1Y2u4UCIuKYmvX5jRYBoyP+S0/fQvdRoozyMjCk4pP07rCalFOqRb
cKrenHRdbMqZWpW6WMiSFGCa0Ljd5eGriyCjL9D/ZC7n966ImJMtZbG1TP1GxRBypKPx40zTFX4Hjf+o38D0MUF5kixZ7NkumvcXcDroRg9Yu0WX7WiEM8XSifi037E/
pRBl5+RKVfQnKHxBRA5E7wnAb4QkreZc8z0CyBkNBKbKiCbRJr2HgYyrX3ljAm2I9eAhsbYpcvuVPp86ImPIqvMW9IDdWP+lp3wSDFpxYxfH9mB4KCH9r+L20vAjqtGI
A/zXER//II61cKZy7W30rsqIJtEmvYeBjKtfeWMCbYjG7kCkze42t6L4BymMXzJtrj7PfyjvZSEse8hkExq/jy57xC4SR/y0U43GFUi4Xj4cxcq5O/PteRywNjFTU4x4
2/bKtlshAIdjfLyduhFtRvJw4gbhafBL5fNcoJ/SiliMqA1COe5MWVNZ1Ccz1aO/pC2WC+rken9jA5fw0Tn6efeX9mZTVH4RJEKx+/iNkdlfxD2QS7EmhakcnXZAOxCH
LTIjStX9R6VDXFFKA2P8dqHQWMcp+nhQy9GEIr+l1cKdG77qT0pL/25BPXQ9DqBy+3l8Tel+k65sY7s/3io4FCAbeiAR+6nF3VmgokG21mQt3muX94/E/KEVrDCktW0Y
WuvHN7HK5u8VzsgzY8/gXrPqzge+g22Bp+dJaQJvBsDz9+N1IQiYxFk+00ZOkx7JX8Q9kEuxJoWpHJ12QDsQhy0yI0rV/UelQ1xRSgNj/HYD2/XI3rOs8DQidP1w+TSY
pC2WC+rken9jA5fw0Tn6eQUsRHmZktzS/wSsNvrSz0eJIeT/M3Zh8N8sd6s8bajzRnXitLBVDSRTDvqWa9Hum5BfoyANlk9H0AVwiMeUB+DawnnXzHJI9WvodRtgwDMF
dd7uNh+twaSOvtD9/bdf9OYb/peoVNvQfZW3r7pKUMZNS2IDPQJ0pY51/+BM3L1NIz5UyXPmhOz0s67qs7RcZtSbGjbPF423ye+SgHMOj4V+OZD3Ub+H/LJDisPmOx0Z
m9M83aNmu2xODXWieni8bB+6rJ7Pt3a6Gzq/szqkCFuRXnhBmcPIgbRkXNDRs8hnc43FJF+BWbFocmwhvA0w5C83/dhOklGBmYexW3sCtfl5t8Ep7g+Bcsa5FBdGc5VJ
yqNkSIE5z+tJl9UkXJ5HT2ePFjGOfzbu/bLM8i364ZqClkFLM0oE1dytpYYlE50nYEpUn23lS21WS4Mj5aQgPhodu8uKySngI9avRWhKPOPOaFQvthdnRbXUnl/SoLNw
DYgdfWCqt/pZjWSLuGPk3gvS5Jzabq3kMreXyEnCHZ90tTeTbQY98sbs2TF733s+iaaZJ/WypPU/tmMJT+68zulztf2KaQyxonKlOtveizsX0+ZiVXfpP8hYjqlIjo9M
S8cfHAMnHvkuQtJHoN6LY5y6//uH7TdgYabESDdmUv9vO2ZHvxsYmSStTH4oYHGPzCc9K5b7KLogASTrh0wjdrWibFDwd//oQsgbSW4OIauawW1RC05RYCd6Kz62gLLO
bztmR78bGJkkrUx+KGBxj6u51cEyX2zqacSqxC4jHYXLg2IDl3BlaLM/5vyHjQNQjkx0LmS7865HLgYNfOOXNO5K8vgG+b08+/NRptxlv5ZTqnLILT4/tErkRWUJKatC
4MgRcgLMHvW1EVwqRkVANTU5YggRLl1M4QIgXnuX59IkkeAzyX911SV0C+IG6thGrFvTQ7UNsu6xZXHZIDyxE/g3PgQawa+i3bftHzua40RlkZzh9oa2lhWVaEAwcfbf
H7qsns+3drobOr+zOqQIWxkNl+0L/TWKqaxTEnfxOFaN6BMLmqonIhqBK7foVfD8FAsCTx46HsSYxXhgFqd5vKCXQT76Go5TFoNBx8QdyrAmafJq4eGXkelH3QjrVvbX
TMLoxSxNOnd/fR21+BrbSBaJIhtIoK/NxPJHpyN3hcnFkimz4w+USi4Lgl7kzbEgZ48WMY5/Nu79sszyLfrhmkbQClGMsJ3g+BoXMRtM1e56fkk7SiK1kYOf6AsKL/ML
b2ArpAJuaRX+Fa12JQSMO131QQRo4WZdw30ciGYxhdFJvm8WBd8Hv9rz3HehZh2g1c8c6POPPDMu6ZrJ+lEdUucHWBvLPS+Bduo37GW8ik+V5uMuBpsZ+uc0zJ+KqbU7
zE8gM3ZxYLlNVA1bEgCizyOq/YU8/cXgQcagjzULNRU+VPq60AVO66vV2HXUQZFp5wdYG8s9L4F26jfsZbyKTwEsB4HzcNO1WcquPm4nImF+OZD3Ub+H/LJDisPmOx0Z
XYUUW7GBEgCVAmbv7f1+FlJuxCwC8h4zEEqpeE5eT8IsBwY3m9/Bjdicp+uaXKDIuEqXLb73emyss6Fu3ZH3p6gD0TwODNjw0RWtcO7+VBf/54o4NnyYxCByEc03U1vh
KhIIpllHS51himFWT0hOCBgxrhTzxczrzaNmHXgEk6AZ9VQz/RQFbvzlGy81m218bgW4MwAQ+veWkvv/cw58PTWuMo4aep2J65DW7O8e1kyzJSDWuFs7buaULdUAJHZv
MhvxpTLGq5kpVRndidEIu+KZJGQRBVNw41k9uiuTkGBJ/z6n9yF58NncS84dYcWmx0TyqlhG2Ef79khCzZ+u4aQxxO9Hrw9C0EaB4wABsuODhaxLfmHk1JAr0sYdXZ8o
qcvCG1vwWhChRX1KPXjMk9xs7oxkFMEOAbaDbVbizFYcDbJPj1mOS19gTHTJ6G6EMEOjQdl0WXupK0iI/UtNszozHfhWsaFQxblnz/x6FPm83XynaXS3vbni++K+5tGw
Gz43xaDZZcXQh6fFntHEOxfDLWnfRQJgQ1rw9iXU0f/xkLxLwK/z6JVyeIhdnuo2+kkBleAQVV+AIbMCZhctjlGiePgGQcx5VH0B3ZnIcZOAPNKa6BhT0CreN0YoDO4K
wcd7G/fTgy41dIlK9oCgPp2sIYePjtYpGvQcdQ/dazFyGhgPXvIqe1rKvl4mTKjbnenH6VRN+bEL9UDc+mWQxAjGKMwsCYG2snvSVYxRLVKfZZUeoDK7T+58fy7SBEQm
Gzt4ryh5/TDwSlb0CrccqAeRYz3m8bvbqntezhFp4UYpd59TSdaKloYYavYbAPJd2URRb3e/0U4myMd2rLFFyD5vroWCASKq7lwmQnT6S2wT8WA8nkIX2iF6pgpHIt3C
sQjgY/a+Odi8GxlHO6sCU/koDsUBgy9mD1XhDE17LQaI/uNW5pfjoVj8HYrM/sGa5duZQYwGslnBemQeQXUPSVzzsg5NyAtJpOhm36VgeNQ7G5YrzTBbHHt3IQRjW58S
lShWgJzQUbnO5j2K35n2mJTPSxQ5OV3pn3j0I3adBYjtRQONL8EJk+0xfNKBowIkYLbGYxA8LBzUqvg7MKc5LhIHQFnorRtiZjBCwHeprEWOMFDvk8QYIBnLjEBA8+5n
bZL3JXZODRM9C97qCB/4H3hRWBBzrmYuy+mv7t7zxs33rUqOOiTSIdhTIMg5HViu0POyg+6mFaQ/GvHYETnt2oplx8KUWpOknMBrGaeLhLv2F6RmcbmR5RMBXx6otA4y
zgY+b8Ry1UBsEUMF7KgmdLg9ZbJU15wVxebIv9bbD2kdnIO/Zsd5fkuA0prnVy+DzFOVgnrx0Ox3Lmp0DOSQWZotM6bgHsnlbpEAa4Y/RpsS8CZBuyBqPRj7gKF6Hoa6
9hmJ3thAVYhFC/hMUUPdDh2cg79mx3l+S4DSmudXL4Ni4uAJpASwBqx6k9cAn0duhkU8vHypGid0vlpu1k8cwncrGYAav0GhVy4+TweBEMGqPaeTmg+W/+48Vght2oF1
qbCoJYej8/r2uz7/R/MSpjLJfXOUgTbqyuTd49QW8PfyCnzYr6/pXQClC2C2PNIHk1JzOCu7Ky8B/Z1CisBzNWHZnAKo5x1ffjYHGWEvqouydSGK7ihlWAs37EGGXflL
UUdzzG0dRVgflrPoGjXBCO4altRaNSEI9X7j395bXoVptieiqqLJ4tCYKHX6Rno07UUDjS/BCZPtMXzSgaMCJCwg23htfcj2PsvUs6Bv2tCRAF8vvEXl+a6Bk4mkHQ3q
KhIIpllHS51himFWT0hOCIkiVs0zQobv54vwyLe9plAsaRbXEiH5KrbmS1mE3N0M5rgSStT4NIeyFQ4Q55W2N2LZKOM2ZudPshAtkn53qBPZFJEYVKbtccWGJl2WYCTt
7h+iHvPT0OAT7oP4QgwHdukPAQRm/I+OqHgpI1VtIKhDzirZU0JeskKO1PiDXSDIdjO2WJlB8bEJfUo7MmTAoB7xMCQh4e+wmDa+78HBWwLemOWIeuk9ccRI1bnjCG21
xT5NSXdcGNZt/UMPvKBCAp0jjdAZzhKTS2EnrwcZrHvZGZdj/+IZlOWJvK/x89hCuu9bgvwv8ZLc0NjXWEfDDEaIwJBS9iBkaLoxewMMrV4znER6bZOorZwgLSb/0P9/
a45AQE+CvRbtELf1zPnpojSyWTM1SY12D//TCzjm4IjEmBPSk0KCZ5KTVBLjAZeB11cc/k0eFMJozDPWYSbXka66Ah2/UNpCgTfNwRS3MUWhDV5ehn/+lVqTOCeMfoVD
YV6Qf9vBGgEN6Q0N2dzSYQt2rGBhVnsmzvtlG6yZzMwcoNKjGDlR74XEZB3rKYlsj7Cv8DeOU27FSDUeWyzcYhCJLOS+HkbD+vejgUAUYcHrYzw/0G1T7MiNZ6XeDLyK
zlA+8mtkzPw9X+RMUIS8bjs+FcowHIPWZY/nMBcBQ16/W52X2SMUNi51jDNuSv8bdJuBBBvZlSde3VhOTgDmf03ficgDsM3KiLrTnZZdw4KTMWYQ64s4weXVnVdlYUv5
5MTHwCPNcns/aMRXjDbE3n33qcyyme/9WmgZIP+ttSRkjb7owkbC60XvVJHOWzyUHx1SI63yOGf2/WKyPz2hnT4jTNY+UwdZJkxFZhFnbTifwqeRVYktIlPugypXTH8d
51fRA18vBBRVtFNg9uvNAS7KX1iQ4axd1RmJT883JxIJDjzjshjuhYL2ARgJPH9ZKsE6J7yHb0q/N+Ch4yIKxrF70n3BsRHmaaeIB1odgNV450IXFFu2+cS5RAcR3cEQ
DQc+C7byNT9EnWoRwp3wjyU46m0G4QKbQhTRTo3VslcLLaCvDmbZLgWeMkrVV6tMWo7ih8ySfZqV8IGhaJyZK+axwYiWEaH935evnpj0ZZTj2KSvYoMebAYY6iiN7r3P
hz44q+lXQItVXdlctRnQN05xGRgOBoBaGvdR/ChxDuG0ouNgomzjPv4xDxjaN1sjF2sY8Vsm7hnn5tNHdKnCsj02+G5gXHeZTLUjRt+gs3z608H93sCE/IVhJUdNWVAF
flMC5EmLGrwW1HuZZmlKNmbqQyFh4PKrAwYYYapM50AgsRUfSt8P0b08j6GvokIyKkHTYLZ3eFVgR6Fcq8b8rN2rei3TTES9zk2nIQf7PAy3i2idn+4+yAXWCD9twfyr
ffCHdPjXseyAf3vwuRYXor7dioBEDdM2Dl9SIooxVQ1xpRpdBfMe+ONT59g6ga3SsXvSfcGxEeZpp4gHWh2A1Z95jUjnmN8ZTBtyiCNYQIIpWSuCX6YdAulibA+DRmmQ
Qh4We3VM1MRqH22ezF6DWo0Vk8xeiKdLLWp3xAJM3PAAqbDTNDlQKl5Kefvb49HCFlm9ghBJpDv0Nii3ZzDQrWdKYeYsrCShEddRIHrerkWKDunv5kxEeELO+mT15JIu
9HG8HfrOzrxBd0aOFH9hLgTz9XwBIedBzYi6EQU+8zp6EwHfuzP+1Br0mSE+tNv7UjV4+ImtmplooE699ttuQ08rAcPbBuITGiuPuutZnl7MB+9cadiOnkTQ0lTocvF6
L+miqaQlfYmU2KJ+fV2uFXyJHMs/fpy1rxbJq97eelGQ3U9q3FAufoBEPwYYR/v1P9TdVdH3dRcn8v3CuUbi6MqIJtEmvYeBjKtfeWMCbYhkDf64sJaYfJwgyF1wKKK3
AiMcNlGgtOiIJ9gdZpQuILYy0QEF6zHy1dQEmi+dH9m+3YqARA3TNg5fUiKKMVUNHs07xlNuhf9xgJMRxSOghylZK4Jfph0C6WJsD4NGaZBJuKkH384qqSJBSaLi/w1T
bZ5ybQCZtbHzpeEJWErnzULX7/adfpk7oUXcyKsp0ck2Z0PazckVFud4E9tsSOAdyogm0Sa9h4GMq195YwJtiOyr55JBhFzsYQfJDhVK9mmxF9VrBh03/w1Eae8X7HcF
sfNTEmierMdVtaQrjn4SiuqJF3Sv01jqk1Dkfc9hiApJtHe3QWtivp/hsvC1hSn2bUpISiB+q3wKiBwm2YQ73MJ4aVU78MKCa/37RhMQ4hPIfPNIrK1HZm2G/2QrQUNF
koRRD7puTVo6QoKmg6rAAR2zut2W+Dx2nMx2gRJ/TVhPTf5K4LWsQm2lY8+2fI8hLVrubUTXMm9NKYcdk65zEvmxsaEZGcSJp23RgRTnZsGjinIdvThfNP7FswxEXTFH
q0tLL6lYMl2Klg7p+E6uw6emElHCcrTqPp5HRIEna4y6zQf1XUajAvWWNfrw8ee8wvr8R9PlYVqzyhPf7vsII16LPD9jk/iKr1mn3ngJj7fw+5kKQ1gTGC/IdWfq6gYd
pYgdozCE/nZqAA5X8w37L1ak27gbfNMn4S4qpSRJCgZNg35foalSW+ooXbW0Wj/uk43gFpEYHdlPhCvT95XSSYieVD2J2h4pFvRXJ1WMLOtqMQgjqX8P8yBGkfqGtA70
8gxgEI+JWHOZLBOcqbLcvuZEx2jSk1AfNAZobBxOpw1r03PWdkO007tHX7mhMB2NO5evjDWEZCRpDiCNJOtYbwF4U8SzUJvUZtP2lXIL23uPnUPjESU2NhaOO/IYMasg
nXUu5tDejCFI3Fncjnlb6c1Tz7YzXkEPtuJnoUccBReHBssJZldH6rHNEv3LWpaCOqhY+iAYqtfAeSj3TO3Avl7c9nxWnMVCweRXox7A/iHWdj0vB9+gxE83j6+UP2C5
eJhaI93iYG2Bs9IIVGqasc4GPm/EctVAbBFDBeyoJnTb+vsM6iswh/o49T8+tZoutSXTutx/XCMOCmUAyY7lcrWPZcud9CPCsYluJnRtIE1bfNxIrGxuIw/xQifpPQMo
+Z/TbLyqBjwBzKrBO9db6/XPUod8eABDwS6yOveSN0F2HOL5EVCOyv7dZgL5vbpXyogm0Sa9h4GMq195YwJtiLj5OK92BrKkaDqBxFKXrnTKiCbRJr2HgYyrX3ljAm2I
nkPELMSQBI3KYVRngPExRm3OxTJfagIEk06Zz4xmxWXKiCbRJr2HgYyrX3ljAm2ImuQH9jq2wxzCfRKQBYDhsTLOmKfN7GxIo0j1RZbbETCeQ8QsxJAEjcphVGeA8TFG
LSWPUGaC1bTTzowrfVxn2sqIJtEmvYeBjKtfeWMCbYiuQbMon/81Xo8wKkuQZKJ9YVhL39P6dNIiPChkpRZQ7Gos8Tt72EqnpAqVoJDI4nlG80tRaBVFIPItqqaQw6EY
WxoVxiDc31LxlrPw2CIZX4dD0yorq7OKRQBnEu3RIpnKiCbRJr2HgYyrX3ljAm2I9rswH5Rl3UkeJz+f63rT7216We2RSN5vQwclLpS7/LqtanQ5QX02hO3/wAtZJz3q
yogm0Sa9h4GMq195YwJtiIPl2yI0B5psbVuXPy4GjxEaQWKbG/hnmtNB3gMZAGpsFpG84WsQo2M2lW8CL7HdIdMxyfjHtym+UTpWsof/Nzf11xD0QHtaBLviL+qEWfQO
2ynaVtTp9nUlJ/kqXE9yisqIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N2awFJ8Z0jw/DBcdKrMh1fZqJ3SiBZNStaEB5FbOxR1/SHPb0iJEA2PI5xU9Kq4nQE
xm3fTEbgdDFOJQM3jQfrLfXgIbG2KXL7lT6fOiJjyKo3cU0ywocpNKp4zXtVHQZKSZXdRwN4saED/s81w/rdTH+zgPoSktDMrJ/QB62SWMMNBz4LtvI1P0SdahHCnfCP
u/cr7V9Xhr0NWCUYNpz7FbrlU7hhcRSdMPTSf7iLd5h+9Yo/eBLElpfqfjnMM+sUpIT4FgSijqNFt69cMXFaC/XgIbG2KXL7lT6fOiJjyKpDk1YGVwUeQ5zlMcyfYXWE
bYVb9qnuR3SJUsMEJ0CklZdBu4o4vmow/uOcZBXUcp9CIf7qwLt9U+/9lG2X0qvjnzkDdlVmwMM8pfVn6MP0k+8qO7Efg8m3NhvLTrNQxI3I/EG6CzJ/7w2hwaqqBDXc
YE7I8HRdiomOjyQ2q1k0NBShIb6dG7tXeI88/Av5bQOxeB1aYBEhpzFZBeNRLDHJVqAzFeXECQd2j1TSNcEE6go8QwXtu5EP5GUZ1WADU425hmMZ5MGoMqgvTRXjzjOw
KRHXipC/uTKgjBnRlOwMkB5r82wbhM/yWqlZiQ5lCHWFNxAS/jZw6A96qepz3j68DbDBZXVA/XYHxKFmuNzdPd5poE47DEfT+hN/h+tRWR2zVn7RDpXjUiQzfTLZd1Ir
W+C5Elv5e65objnGA3sRO/w07NvtuqNA2rPAF11UX9admhbP8ulVJoD0NTG1OWEZNpTzaST8AOEDh8vNYaPJFZHbJ51Mh53PFBDlHP+czmJW5EPzpagrDRGy6BushIDu
pgXtC7GQUd8RP9PCHpwYBwCdOaNWWhjT13QwyMixRZmuHm2HJbKRjsY4/1WcRdW3nzwvUjsEpzO6IAb1jllp3NhiNQzYvuy4sVLxmegsB8d78PjIYfo1Py8RU7HKBEHL
nVIicgV0AwiKaOWZEHfVUi7TGzTJE5a3J0MaqQCnavO7QYp2Pv+BOtYgsSDDBtNqCLAghKA2YaDVmvzKJLvAnVwyIZJgolqJEylinDKkvNSslUymHmIP2oMC6aOFQbjZ
gq8zCNh4hJeF3T1jKWc9AYYABjm14gAcho91quNd5vc+0ltDXCvh5L2UJU8oRheiAJ05o1ZaGNPXdDDIyLFFmSka3cK0Mk2lCgA0U+EQ55XV2Qr+Kpi+6S7g7Vi1SXBQ
/b/oFNLlWrujL8au0xGVPjPOUwJ2jvs8BlP5P+jNDe9Yry+5J1SUp0Wrrw9eiBps47oGd9KUP/YQ0OuEl5zGRWQF/z46i85RppQFhS6Z/yvFD4U2EY+RwCG0ZuZMLYF4
9H5ojxdoFGD1KvFEAHlVCMkFuEdor1mp8IN82deyT7+NJKnGePQL8k/ZCy4im+m9S6XhH46R7YF9vj8zSKNQX8p8MzZymID8RZcLzQN5g4K/ZmatZ8ol9dL39Yz/5ib2
TgcGvJhD5IQo4hk9XQKZSepuNQBkJGIOvHhYkPCY/0WSaJeCYGYIMsZrVyCPLMIXbCn4ciGSyWhk7pd1M8siQ0lQ1knTtBtp+rYDR9CWdKQFWoZYE1SKLIj7KPg34548
nER/KIg1OMaNdNdyxVjBZ0REIBBTfr02frbp1OFM4TgQLsVeD52bCwE4xlGFrvd/ecN0mDlyefLoZXGmNw5ulc15In3Rv3xIJGDSEqlMrMbwIxs9btbSw2+xLYfuXy8T
7xmOVlHAxOQo/NV8oYNNSCD8xQp5q5HU3YEQKVZYAJBslIPfSx+/ru+b01000L0cCGP2siGdqzWVmsPaTOVdp5gjYRvmgbkyLZF3TID41An9lQMvihlcA2gqxa4WcZjL
5k6uaIiXJPmHZnuaUVNcZUjohphOh7YqXYtH+RF5EfYK7V+EbIcdo4fqBIdRknmjnxt+kjp9q8gLW4rSNLJNxlUDyMhUVkRU7qCke/vgTFVkLIi5Ulhev3WM1si8dtXu
v1jDYKw/TXJoKlG8Lm24ecZHd5fkn9OtMEPZFSEuT+9aazF7pf1YNVA+IeOQZ7ieZlYacA2md3AHY80/MSsZU5zSftQbpECHUj7OzOrkFhsFEVeQL/m8G4HOHROk1Jza
ejhiv58R+liJWql2WYWmT/ya/D93nkwfCcsw+NpenYdM3W/Hgp4CNIheFdvYlDiDE/M8usAQCAzq384FqnEgSdocyJxjX1TV55j4L9vXpUO8MV1BhzpwDIQYbpFg0S6y
PtixNPPazkOsFbQPrrwE0Durroazy6tz1E0bzTVX2FWrwGUSxegRQ1UvbCoB02Sw8j4L+7tExny7xz6Adc7+dBWTn2YknC8s6kylDm3b+6Pp4qQBo7erK3viC+Fxjs6L
SCn4iJflktWW2SCvT5PFJQfJUWQaHgbFmYkzumy43DLNFVwP0H7DLge7nHgP2+ho5tyPVZB1QBh0VaWCiVXucfsSxJjuG7olHOK5SW6VL6jxUEsXz8GyUTJuzajC9ZqX
iTAjpYz8Nm5rjB5vyb0aUPFQSxfPwbJRMm7NqML1mpdhmnZyfyoh9+BuiQCRtQDDnhvyxUlkZzI7mfkCyXeJuLBKhq+RcDc4dlUb+zh5sJsTnWYbC/5NeNLyOjNfTDRb
KsU/sOkTInMGJ3V2ccXX7rk3dppmklPh6m0LZQWc51/wXJCXFhEbc7Qm0VA8wIdMsFMy/PAkwel+Myc6q802RIrTnqKgSMG4/WdJ5306z0/ZiD9hEquIhvG4ElZjBc0N
lM9LFDk5XemfePQjdp0FiFl0FcKzx0/8nehGztSzdV9UAQ0HoJTtw8EBbvYXQeW1nhoFrNIoRz+h4iJa092utTISIfDYraKBv0++ANpxrwedG77qT0pL/25BPXQ9DqBy
zmhHYjYrWLLO5EHpZPREXuaM0OOLmZJyelyoqHiumW7bhY6dYEMa9WZFvke5Epk5kFCI9Fy41UYrKg2BK2xWNw2Nhf3/DT9SvpeGDtAUlUa0iHIiCEXxPQtEpptUQILy
hppegyGEamTjAv7TCz8KIEm4qQffziqpIkFJouL/DVMmmRPqUNr4gHOV1GTe40ZZMpUjjQ60V2nXkY5MN247kSJC/pHPWY41zPXs9WlgeccTD2iyFGznju2Qy2IBIRwb
QUcZv1QyOtyMsWATDVgVo8iQOPuBO1doWDVVjVQdWXVYomWlYDItXkQNuNMiL2/w3lzzL2RDiyKRnUClU+XbghDnK+d7Yb7WjbVt0UrEEp/3rUqOOiTSIdhTIMg5HViu
mj79Kl4pw92HI/nqwRXq0S5ADKsw8QqgNQWmfh0+lm25N3aaZpJT4eptC2UFnOdftIhyIghF8T0LRKabVECC8t8olKugEj5p/27WYroKmfNqLPU8dD2yyXeWsP7Ym2+Z
Y0Ld4Ou2cLddGwXnv5hcbJENZxjS7cL0lEo7FE5arWtD/f+lw65YMQQLi35ybEutm9gTYeeU0JPm/IMCBezRabipdSo/aOPVGl8a9c7UCRwn7fJ486C2XyZI1RANxlKK
HQ87wozU++4tjaY5ADzpvJmW5losEc1LS56ZJFZp8xwAPM4tEjK7iYsN5uMLgI38KFkwvztUhxnKV4xrbcYlY0R4YPV7fXRdo9Z2s8VDdHqS66GGriZVbWQMaHq1QE3H
OHEXpDUYnvEfK2C9z3ASn2LFziol+uXDe08CsSndPl87PhXKMByD1mWP5zAXAUNe5riNLq0vRi45TLchusRZx5IiuX83Bbgp0Z7pCdDWToprjkBAT4K9Fu0Qt/XM+emi
d3ZVX5LDasvXFGwOrgHeY3SbgQQb2ZUnXt1YTk4A5n/UIbfQtzPqFmTT1d+Jk2i/U5sfrIsuBQu+vYP36m19UHTnVJGy50OAZciu+M1QcaFlG3HCbQDo326xFDzaMCmd
EIks5L4eRsP696OBQBRhwckVPabpqij0fTXCtJF3dZKBxhWz5iI4VItjYwTATDBX3vc9aqxMGeFpaENZyuJ9gPisO6YsUXmnG0ewLY15Ny6bzbVG5eG1OPKVux52oHnG
nWN17tzWfU/U2AIe1shYUUVWK79c+NiZAjTQZqnI9IEf79OYg7PFprzwNtAyxS8MMZ9hDO6WsKPe4PgILIKy3YQjaKVixVRzWt7dKkp6r+10m4EEG9mVJ17dWE5OAOZ/
Hti6DiccUPFrYhwhdQMP+Mrfzp2LFqEYzIW14ZHqeXXkxMfAI81yez9oxFeMNsTeZ8OAzAWleVGyA0HbOJJtwnSbgQQb2ZUnXt1YTk4A5n/FlNBVTq1t1DJrnkikOU+X
vWRUKqVhFhkLTv/mXkgUTtHlKFEiX3hS8GwLUzkUmckpq7c9DrjNbfsn1mofbMFQsXvSfcGxEeZpp4gHWh2A1QJQ7Md25wSmVgAjGZN9N66fwqeRVYktIlPugypXTH8d
aZjTs6fKXwT6FWsJQE7Kv+0vQPlw3BCax9EpEtjnss9Eq1C1+b7qMK8et+yzMDA7T0hr39G6C7Nbl72rjFiM4k4HBryYQ+SEKOIZPV0CmUkoMDjK9tC/6sbAA8Ikc6YD
zl5tkFu+up7dMUFei2iioilwUS00x/xiMr5rzrp/6CQx+ZL8Tvn6Lx5iA+ROuEXOwnhpVTvwwoJr/ftGExDiEzRuBEbXQnBDO67jpqHI1/QJ4UVjc1747yrPodKjYg49
8IsmV1cYs1VOKE8fMtOm1vek9PVWdF+tc8dMYaYO1mEysJ25GTPKWsu5Kgw5yOCnI9LRevI676yIBdyEQzCeIAoMtDSpAI2i9S57Ej8nIHmznSBxJ8oBYzj2UQGnCWzX
CM2PFlJsMuRYhivYT8LyOLkGm1zFvD2MnrBxz4gMb20pes2SdP1WuTCoFV1S3eMGKkHTYLZ3eFVgR6Fcq8b8rMnUxnGnfX3ROQz2rKFZboi3i2idn+4+yAXWCD9twfyr
ffCHdPjXseyAf3vwuRYXor7dioBEDdM2Dl9SIooxVQ1xpRpdBfMe+ONT59g6ga3SsXvSfcGxEeZpp4gHWh2A1Z95jUjnmN8ZTBtyiCNYQIIpWSuCX6YdAulibA+DRmmQ
Qh4We3VM1MRqH22ezF6DWo0Vk8xeiKdLLWp3xAJM3PAAqbDTNDlQKl5Kefvb49HCFlm9ghBJpDv0Nii3ZzDQrWdKYeYsrCShEddRIHrerkWKDunv5kxEeELO+mT15JIu
9HG8HfrOzrxBd0aOFH9hLgTz9XwBIedBzYi6EQU+8zp6EwHfuzP+1Br0mSE+tNv7UjV4+ImtmplooE699ttuQ08rAcPbBuITGiuPuutZnl7MB+9cadiOnkTQ0lTocvF6
L+miqaQlfYmU2KJ+fV2uFXyJHMs/fpy1rxbJq97eelGQ3U9q3FAufoBEPwYYR/v1P9TdVdH3dRcn8v3CuUbi6MqIJtEmvYeBjKtfeWMCbYhkDf64sJaYfJwgyF1wKKK3
AiMcNlGgtOiIJ9gdZpQuILYy0QEF6zHy1dQEmi+dH9m+3YqARA3TNg5fUiKKMVUNHs07xlNuhf9xgJMRxSOghylZK4Jfph0C6WJsD4NGaZBJuKkH384qqSJBSaLi/w1T
bZ5ybQCZtbHzpeEJWErnzULX7/adfpk7oUXcyKsp0ck2Z0PazckVFud4E9tsSOAdyogm0Sa9h4GMq195YwJtiOyr55JBhFzsYQfJDhVK9mmxF9VrBh03/w1Eae8X7HcF
sfNTEmierMdVtaQrjn4SiqYBhiQ8UxtI4ot84xQ4ZLZJtHe3QWtivp/hsvC1hSn2bUpISiB+q3wKiBwm2YQ73MJ4aVU78MKCa/37RhMQ4hPIfPNIrK1HZm2G/2QrQUNF
koRRD7puTVo6QoKmg6rAAR2zut2W+Dx2nMx2gRJ/TVhPTf5K4LWsQm2lY8+2fI8hqrL5Un/9g10HkBJHfwNV7LEfMKFG81dbgoWa3cWIRj0V0lxjabrffIfqwTcuadiW
SLjQLBK4VSuJ50X21lZfm2isBGO8/WMYCs2JEMZacgkKdz4BEYw1NEcL/SraV3IqX+mJEErLd3uiwtIPgw7x0l0KzcZ5vDEI4aVb/tz1rBw4VaP8oshd06oqOqEc+8/C
KUEZj6kcilteQwVS109bZWq59BWLxw0XA/yVEn6EmmbyXS82dwpXUvbiihaNvYnLlo3Yzx4EdJM2PuT+4xxyvMxdMtNEO8+dMBKo6z+YN7pumUbSf0O9UIUZpSOoUSy3
Xis/S4KN6Ar4m+1jxKk4gF22jxj0CEI7goXcCgkd9jx/TnYnnXgsJrQgXYcO6t0qJm/Zw1Qp7wKQG1db6frVZwDj+hZBGw4kuDDVZd3K/mPW+yKi2ytmmxPvDOakqR2H
2ZkZjVZ7kUZAEkg4EuVt8oY2A/SPw17VI2pTLs6OOSAUcb771VSXb59d8uFE8fnFTgbvIsNibcIQHrNIz4tJPWyfK0/yMkGkY9Q91jhya8TvXtARhnKKUMfMhxDHzkUs
zj/lZ1jbQMwp/+TEIv2qEC9VhLaLmclfugonzEopARqWnTJr/9PfS2jsaIIAZ93Vj51D4xElNjYWjjvyGDGrIJ11LubQ3owhSNxZ3I55W+mMSMKrMfEM+6tJGYrADkgk
EDrKauVyOeU8+13wOug5vJbv+dtgp6ZyagU1f8v4Ajkm0FHyfdi+bMxGODjau9D43RptSD+5noE+1O+6vxn3sHjnQhcUW7b5xLlEBxHdwRCS/5ywCSLuhYTCoqQH5eFW
/UiTKUJyKWv858XQ7e0SSVxlFOCczmV8mfE+Yq6yRVwyzpinzexsSKNI9UWW2xEwyogm0Sa9h4GMq195YwJtiA/hEA/xXAycN1N4kxQDTUJo/Q7kxyeJZ0g98WS4h+s7
JcXG3xJ0ywc3JUU8EJSDCPEvm7a+A73mHkS/xwmD5E5PQB1KjT4ijF3ek5qmB5wxkAhEfXZlVZ/3y6utN9jMiSFf2ns0JYHzzaZnK+qEQzSPl+50Mo8zL3aZf45h5nFB
TgcGvJhD5IQo4hk9XQKZSVhf2ZOZG1Nkb0FUCrDRxUsJ35iUWhwDqcmI3TqxXSYPX98BFzhAJ6GteaxsTUwvs/DxPR33mpkusJbQM4SIMVBPQB1KjT4ijF3ek5qmB5wx
ZxyZQKcsjlW/ZaKk1Z388bD/xX9HeIOJw+G0usvRGf4yQgjiUKp6FoDM1XkQXp5Qyogm0Sa9h4GMq195YwJtiLDsgheWy3/kN0E9WMRXgFew5nkhEoq3RLbFQvAcS0bU
FpG84WsQo2M2lW8CL7HdIdMxyfjHtym+UTpWsof/Nzf11xD0QHtaBLviL+qEWfQOfO4eF8Y/ccO3vBQ+dwrM9249yqOPgox/MoPbrhsZmZ1PQB1KjT4ijF3ek5qmB5wx
kAhEfXZlVZ/3y6utN9jMiQD54SpDMJany4yrHdc5gAryhjF/PUd2GtgLvzbsm8P28S+btr4DveYeRL/HCYPkTk9AHUqNPiKMXd6TmqYHnDGQCER9dmVVn/fLq6032MyJ
IV/aezQlgfPNpmcr6oRDNPKGMX89R3Ya2Au/Nuybw/bgz2bjvXY5Jd+Swcl1AIPS6HETvUzLD6dWvhXpMplKuAby2vpc1iIU3eKsbG/msDUGgyIc/DkbJJinnUgBuzjB
xFIiWVe/4Y+abJ1ziL1aRsqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iq8xb0gN1Y/6WnfBIMWnFjF8f2YHgoIf2v4vbS8COq0YgD/NcRH/8gjrVwpnLtbfSu
fXwI1US6C8zsPgh8VL6iqwmbzPExbhQpAgTRi/SqjyCFOOfMHFqfaeqJo6u2eQ3aOEvXZ1O5PV8FmZ7CoIB+5YOSgFVp52grd8b8YQv1rOHdco7jc1bkEnmGPw8VLPgD
oLLkqzo80iqutKG/oMm45S69oAt7g9muyBHm5/StP8F8IazR7hS5Q/kN2j4MNXl9QkmDWdh1JDYfrPZYG7a/g6N2Rux0eMuqRWuJkRgMmz7Tf8N/Zo5VyS/L8qy2dSyR
9DDNJx/NPKmBBKyXzOaVKG2bOp+4jAYI1smmPcfIss5pNgHO16bT9hus2RhFPNB2/zmHHpiv6FmwCd4m3PY6d4pURn7IHuTgGuCGBFBUV42lFl7jBBPfwnizd353maA8
2PSBwYVp1vlzrCmOX03XoosLM3CUR3F2R2uWU5OPc6gsn/ygA/vknaTcX3z9qvOUjOjv+hyOzUNSI5pru/89MWuA3iODO5dbWkmSW+92vQf7wdI5B4HzJ9GN+J2Bg8PZ
8Pf2GGiWE6umBBVdXWgOqhJb07ktNSo4Rf0BIw+09qT123y57EG8ae3hAx3zp+HXiO9746WZsEhOhgTCAikSQX4pzDiGULvlT+rtiDYII3oC6MZJFXdzeob26QyGg4av
3AlwqB9zDYXdpzW2MiLoz8vznKRQlXSrvSqGFAIe7hViCM/j1ardUdo07iatGBM/gr6Kc7fX7iB2d8iK0NRdYKKFF9Apo0OUW0rCFhSVBGlUUYCCDUKG2ZOSWJ/MRVmD
f/V66gKz9EswhH1EU6icXyglAUu0zv4oUT4DtttXZ3jruMUzRN1pxjW7m8lkeofwYGzED3ftmwVbCBy5/2d1/gmSsEbth9ofOsqN4RBP3LvjePhnMpjfx2t4NToKtJCG
qPwmw6zggUBJHzCWILIJnQRofaOZkRe4j/7tr/w7ModHg0X+2F88xJk4mZkerlB/dkelbi/eD7CZzNekeXTDNkckUUpJmX8dt8H32bICmuEiNq0Ea+CV0lIdKhoPys5S
RQtq0j0EM70wMLD0lNFgln/0M4ImSnJM2Im/MPFffnSaEzNfVVANeg90trISwHwT3kPHDNyvoGT+wG9FmHcjNAC4Q1tRVaGZQZmrwRo6c6ARyWQDtO5Ej3oaawJqGm/r
zUIKZJohsJfjQ8SK5hOIT+1zIgJ7L2c+1XW1dJh1/t210jcgq/gthtIlUQGrdaQFhfOp3YUbq+6JyOgg8mJ8IfWJ8t/ek/hhBivLpUS+vSKuKDbCpBTxEJHWohDZovv9
HqGS190AW1b++SxgVVyX0ihaZC+Hf5vPsSGp1R/1/HHhWJ61y5hGMwMuRSUBsFDE/rNLkp+UPBt2nSClE9SDVf2ttEFN6Yj0m3P/NiCnW/domIk9fUULu6HunHzQ814x
HkqUZdGHJ5zoeK7Q3gVMVukkVidbj2/ubMkIcj3FU/yKqmZmaK8Kv9MtD4Wi/53ChHKc/+QOWLnuVE8PeYfAGM02vFyLPmFSFnMEhTYoGTC97b/Gb76reooYcv+bmXRj
r5q0X6d5682A4jFms8o5+50c5qSAO8cNgmEoMU7Qxfj6Ca0s2TskbA+ryslzmxxeU6AiQfWj2X2e0IzywvCikD4ble5l2X5dov/VQTwAXj6VW+d2BYLnc5gXogtrOdy5
ynwzNnKYgPxFlwvNA3mDghfOktSGw/4kBrr5n9vZxRp2/Its5fXX4tfPt/cl0mzZU6AiQfWj2X2e0IzywvCikNHzAbo/rhXpFBTDxgDRqpwZlOQTiijDUBffYYf8U10z
SVDWSdO0G2n6tgNH0JZ0pBr2xtmQI57JcPIRDcre7zRw57HiY0LhdQJ6weCykjNDTQ7lxUwYiF8hwLJvmiKlYULXpA3cTTK/yzuDMBkSYSnKfDM2cpiA/EWXC80DeYOC
RQP48pY64+WHHK/DGusj+Ro8LvobPKKeZ7KC+yZLlcMccDIdrylebhVc/TPFZEV2HIfIoroVeQYaAxh6+xC9IrhE9tyRnA7I0v1JBTwq5qB8ZTrukTgobwHfpiU+VzAK
a/W8MbJyrVylN7k8P/436xeJC7A1Q3W54Sl5N6zoD2Grrv7ANdeIticFFzDzyqhb1M8juHMoMRP7MRIVIYpM3cMwQgHUIXEIaazKA2WXf14T8WA8nkIX2iF6pgpHIt3C
fd/QLxQdjFA49yqbBVAEZvc/4o441DuHlZO0rOkj3hx939AvFB2MUDj3KpsFUARmxJlBz5qjfjqoEmx/3dv2O4q763yxtgAMa5rd7Me+ez38mrKLBBOc8hiV5jkEd0iZ
C9AjIg1hNV6KBqNqZrJeYEfoi0oZDEvHEQYZ/iidtp7b9sq2WyEAh2N8vJ26EW1GTMOhBksEz9x6pscMwVmFyx92bBPgXOJWkLB4EEpEJ5TrLQkiEU6/9bQETXvxoY3p
WzxpfbAEPk4jrAK8arpnuMVJ3YuiznLBoAZ/M5J17x8pUzUhPZeVC2l92u8lZ2g2KWewoUTksIi+/LfLJe8qf+Wd3Blv9kScGut0wciO94QWAZQwBvsebt7ivmZAMm4h
BUsdlkP5SAKfpZMCzoYQyAIfze/Ff9BY2r//Zys3SKcyhlaQEubuEsz2BHCFsQfDw5812xJ4cjOxiHkn11KsmKi/MoWY3jTzg3ReY08cYjSE0Q5u6Nhnf2QztZsgunQB
dbBPWhrubPpEamW5ktjxtHBZpUAwwVo7Eb9RQqS8KXqSccxXKLndRIf+wYOmeAOknhvyxUlkZzI7mfkCyXeJuLBKhq+RcDc4dlUb+zh5sJt3cto8Oj5fwYtwwBrOaD8A
KZn9Gr7GrwYKd4z8zLOLtOEVeYBtHot7eYFbO3lBiAFJuKkH384qqSJBSaLi/w1TpuBHt7bwxmfEpC22uDLbcLjxuHmpe2J898pAmPjUkjzHClAkSzOWOzwCRBY576ei
IkL+kc9ZjjXM9ez1aWB5xxMPaLIUbOeO7ZDLYgEhHBtBRxm/VDI63IyxYBMNWBWjyJA4+4E7V2hYNVWNVB1ZdaYPzns1JWz+zlBHo66WNPvXOtSUik6R6ZWxpR2B8SVG
4BXXffItfpenlpC7GzKbaI7XVL0ze9KBxGHhzoIbtSOMMoiGf8mUk3RQMKBBh17PW92S/5HbSxmJC3pBVA16dh0PO8KM1PvuLY2mOQA86bxU/mKQpg2+bFfKdG2WgWlT
T6Z/ZeQMOGgudhSLEaTWChxTFVy5BPwSqPNEZHPxKbo1rStEI8q7M2V5bvAHWK6nhaY1QlSw67NwJWVP4ff0nSIHTB/lhWIExAPxQR2aMt0H39EmOMVMnxKb/oAbdJxx
qzPvag2JCprY9ytPrR74OhCHZNzAVf3X5POHCF+Z30Cb2BNh55TQk+b8gwIF7NFpgyv7o61eEelGae8VJTr6UNxhRwU1KPtb4NXoWLjVHq50m4EEG9mVJ17dWE5OAOZ/
VcLB0nQQi5+zTFpI2x/zwDZ8cw9UDaJHUcgHOisFONFvZz8WHCAWbvpxrKsuEkA/5Z2OOsvnkjWStH6RLA9c7qlbujJ2gQjMrLlvPmxd9rTXGC1UHnqfR1rrqc92yyvU
md1fvQ0NPO48yXTcBWtt8ikINysCNi2aVp7J9/SQ+vw1H8zM1uO6YvbUg1R28o9RbNTyQhdZ2hWpO0d+bXeYD7nQgsk+5onzGLGJirzVHpDlR1U+vVS61CjNc3PTG92s
UOFJwZAyKwEwZu7HtI6lfMeiKBzUSyOwsHuFXiuO+eZiLeyb8ViQs4vr4f19RSjDZOfDb0YOZlyjO4u7mVZnNuskjn05q8qJ3s2qtunTtHyzq8pJCQ2z4wsUah7duTKc
1LO1RcjTCGYbv33V3bkMJRsLaQnWxHP8gWBecSwi/AoTMC0wydqZaECpt0mvbtFZoVUg6+gcBFVkYyJJXiA6R/1ehELn7n3el1rN+ON1E+b4n2H4qi8YEwJhBr8yPk73
2YkfHBgv3nEiqcvtUg4ojFgF9GkqvI3T532KH4N1qB3L78oFxG/Lp76qf+XkryUKdT25aw0JfFA6cidluytw5R0PO8KM1PvuLY2mOQA86bzPqFg7FhmREWDImtxIbEU6
DaCxRn5y2rEHEv9pMyZqi7a3169EtIj5unZk0RPZuS4vzxrf/MDwr4sEqx3RDrfL3W7CXfAnjRNyYoElAvGip6ol+O0kPoJfYtPzqO/zqZmYni4fVWa4UMaXa60Sr71B
mwuXfqGB6cWmG+FjWgFOm8WZLGoQT0X+Jkw7ifGsGaFO9vJFHme7Ip/aFiyFRb5T5RoVl7KaCH1+jl4eIC+Bdo8FiCIckupGEtCTzEvOH3HULm1oaon+S5vC1scfGIih
Hi2Fm3Qlb3U0VoE5Fs3EypIcVks1njVExZropNmDUNfhN0kcJgoxJamwDzJ+PVdY3tg36JZIjTN8D7VQ9R/Vsk6HNjmcMIvy9yYWlRSw2RxZGWCdjV1lTF9PcKCeA6qE
b5k2sGuzbUnpJOskFafGephtCRQyiTjTV3zubrbSyYpebJ+lz3gZ4J61woMiX9PpoT1n22ukde/n/K69KZKPsic9TI8VVfxwqk77JJv5rcibe6h1/VxL0rZJ3K1/yYgm
KgwIUH6iejjq/p59X7pl/czA3D1Zbfj4BS1MRab1+jhYeQKSUOmOjQ+Zx9etXQDdkN1PatxQLn6ARD8GGEf79Sceh/Ex52ld6mOda6JoRbrKiCbRJr2HgYyrX3ljAm2I
LHI6DQTLtQi7aiPKhw8s+QcmXupvIc4qQoymKMbXYJf3TsgmpCGrpysRXSMwFpAAZ0ph5iysJKER11Eget6uRUxUFaKX4ggdIV7RqN0owhq/dk+zJVtJMN1i2MInnzXJ
2EXKyWM0Qh4rCLYhalHQbDKwnbkZM8pay7kqDDnI4KcfLzNinDhcf/aK/srtlz+t4fdACgs+DxdUuLRwJ+WQs4OwNrSrtilKjVU/gkbmIUTRnbEby0nHesC7ddwZUMdq
MrCduRkzylrLuSoMOcjgpwGbagVpe5EfgSgqgQZ87IuBGMEp09+885HqV9v2BVQakZbs44crzKsiwk+wf67VJ4dYUNn40WY/ypK1Z0D9fcPj2KSvYoMebAYY6iiN7r3P
OUJ/5IpCbCI7vdxV97PqkmyR406TEovbyvI+VhDEMMetlj5d1KQfiVjqiZJJY1NXZ1aMaLvyJ2hb25eFtUuNP8wH71xp2I6eRNDSVOhy8XqpohjaHq1xXJtlIoaHqC54
IKjL/p24Gbb2kM7hCjzCmoTubAX32UJqMPz+p5vmoX+Bev9gWas7Eq5kZhu4nv+nMhDTuPSCqOZoNrYmNBjl4b92T7MlW0kw3WLYwiefNcnmAX7Z22BPts5MH5ZFO0wo
sqpEC3VOyOzLP4D+U6xlGjPgyXg7ZOcU9dRywCHIFZ41/VBz6HmRg8mLB6sTNbpgrsgnB9zSjYueDo1mIF04OV90nFL5uPWxM5G4D9e6Wnexe9J9wbER5mmniAdaHYDV
N9vpW2hd7NSCbsU1vShy/aUmJYOGfyW69NHhdKdtiasqQdNgtnd4VWBHoVyrxvysR9rOMyldYtNAB7cWVzRcKN7YN+iWSI0zfA+1UPUf1bKq1ZzMI/Zob+dgiIqN8VcD
HmcEzAtP6wSVwuUCrOrzcCHFvNiqQi1T5MnwKL4z2nLDyVPFyT9mkESy/hN/zYLAzmx9ZIRnJTi2T0FOnSxsGvmxsaEZGcSJp23RgRTnZsGjinIdvThfNP7FswxEXTFH
q0tLL6lYMl2Klg7p+E6uw6emElHCcrTqPp5HRIEna4y6zQf1XUajAvWWNfrw8ee8wvr8R9PlYVqzyhPf7vsII16LPD9jk/iKr1mn3ngJj7fw+5kKQ1gTGC/IdWfq6gYd
pYgdozCE/nZqAA5X8w37L1ak27gbfNMn4S4qpSRJCgZNg35foalSW+ooXbW0Wj/uk43gFpEYHdlPhCvT95XSSYieVD2J2h4pFvRXJ1WMLOtqMQgjqX8P8yBGkfqGtA70
2JJ3Sk8fb1/yhcNU0fatv8sUcoUQdTLLin4fVY9Jxyp7ugY0+cVDMdTs+1+j7A8FXuGvuQfsUA/TbJIaMCXnLHANUkp5GfpMLoRUdsJuldL2Ic+rvQHDL1qbQbCdq5+U
bJhJ7g7lXPQmAxTffeqh5uVls9KeSGHFENkljzg5PuFis4FUpvgZgkwYO1vdQm7+pxXA59ewkEz8gMhPjsSHT4lnRGsRUtiHFsgFGGlZISCjp4AQXNc8zVTY4BwW47Xe
J47pl2ML0XStP03yW+n5ScYWtswNbeKOoeBtvYv8TsDRrTeHIivPGLIN+PUq3g7LuUmf74jaevfgJQPE3/ftu0Kv41QZo6XSTBJVr8DbY7XsG7AJfZXrq3bYzxgBw1cj
Cxvo3QRyv4Ovwj1JdHqUsP970MMqfDIrerwDWztThabwMko2/CtY06emUHdvU2hSB563G7mSsO3bx1zdILgFQ8AVb1B52I+P2UXOcAb/XRX2HuJhLKHqVpVDRXVhL6V9
pQqjkG+2kViz6WahSh8fp/Kzl8WGltUIPrZVc1tD0O5VEBIaCtte3TuscMd/vtsJjjTv75tBkigkmUFCvXaLG8qIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOej
8/I92qitxsDg6kcOMEt5PZERLsC1IlWRGd1c2zLeDPaxH15cFOQLBIWIiH+WGMx+bj3Ko4+CjH8yg9uuGxmZnYEayJwYGQ9fRzfY+QWc56NPEm5M0bNbei+lIHJ3jz7J
kREuwLUiVZEZ3VzbMt4M9p3uOwBJwVD7uk9dc5ViOBNIfJLwI30qbKjuXz685Hs/2oRyWKk0HGc9kFJ1BBrZD8QAKP4QwhReDUPsoxit9UEMt9N+4L5xLHYVPmSHgFqN
5BwJ5r0dhNW6F6o/grdZacqIJtEmvYeBjKtfeWMCbYh5H24Cihayu6ZOI1RLHJB7+oI/4T1qcyUjIGdq76uadTZxRT+N0mEAyoqxu7WaoT7eBEehDRu5tBQw9W4ARUw6
m/9fZuZTcqe2QwbCO4TAXo3gXKnAotmwW1c5LhsWjsySHFZLNZ41RMWa6KTZg1DXAiOm21KkMwRljQR2a+zbcQQTrySqLEIU5UWkLUj3hBRx4YFCXlZhL6e6FEZpvg+L
yogm0Sa9h4GMq195YwJtiPXgIbG2KXL7lT6fOiJjyKrZ4ISu2pdxquoXYZCAXRebSZXdRwN4saED/s81w/rdTK4FkAYo3yHGM9VbVO7jEMpUxpQyd0HAX6TAySxe+F5G
oFN7gHeT+ZseMhR+qjrtIjurdLcxHYB/lZFOueX3H8XlZj0SNRUzM3DQ8ZuBA0al3kPHDNyvoGT+wG9FmHcjNH+3hIdGtipNIiuT2muKQsjOy2E/N/5dgn3+aMiPSCQI
1qPnPPeYfU5BZWGX+NMbPYnzke01u0flDLNsLDGpUvJNrOe0POlmnvEHzG3DuAc+oFN7gHeT+ZseMhR+qjrtIoFnzr/WoRymbkMJlikvBBGHJ2By31M7eIPw/khJQNBK
s/VBL40KGn/lFEimoHbsMJQcVJWN3VgEeoqzEzbIFtEfQUWHnugczoSyzunTWg8Oi2UbkTDSQSLUdRI0WfpqZLiqtBkNzBa6MNy7BH4VShVr1LaucHL4cS5t/U1e3XXA
jE0gLrxxSiQHGOuruf9+W/YSnlaROAucQebMTRh3qXv6HWOui+a0GxjI6j2GK/X8j4a9Ox8L6YGbyCIO+vFiV+4AsjgjTkYPVw4fWswrKBE8nmzFBW7W1vl11zaYnaq+
vNccan9pcYiqN7eyQDfqwSZTO3YrelFdHh2u/iLrzai4bXgsybWK9RgA1+aPyZVW4M9m4712OSXfksHJdQCD0pFSkZ0+5eQqSO8On0Ga+7V2dvXMGjwVXjCUg/p5pJ4X
tAx/7Fck2HSvr2qkIzvE0cbUhHIkX8N8c+X2L1nCNNmCrzMI2HiEl4XdPWMpZz0BPmFa/WiC3/MZJxgu+4tLlooO6e/mTER4Qs76ZPXkki5bimKLye6bnHi9nsmi2Qlo
4tBH7zqRCJ/QOYX6yL7qRqzovax/m7pfoZo1Add6OzzFo/JgoBVrzgtqJK2G/1Dn4wRysSxVZIXUrujO7Jd7koe5WxplJU2fHB6zCPkQPKGCrzMI2HiEl4XdPWMpZz0B
wFG4Be8Ebxr5mMQAQGXrAmOk7u/mZAKfviGWZRMGiqVB9fc5ozC7fnp+vT8GaP3CuDxrCNGZHPlVNcFhFp3x4RbCyzTrwNo45yVuASJW5eYAnTmjVloY09d0MMjIsUWZ
FEFvQFYjh8HQxDHv/3OZGSg+h+K+mff80TFqlEZdqMK48C5vmCBZJBn4t2/VsmqnZHgKd+3gNjeeP5glZRtRdSr/+4XSbEHdAYME0wODjwLsC3LNDM28sRNYL3lMt1cg
UxTd3j1QT61TqG7IDLBmtYelvnSUqKGtzFvdIIEOn08/ncdS4Mnht2/JnTbF0tpjVIGfK27lp73I2GRoZTk2Oeaq6TAXQewkxoKIqtz2Wm2A2jDwFRxXML/sMEOqoy+s
ClWnSBAGp+eULqkkPNAj5PaYsIGffv5N8A8q40a1fNRo7sgOvdglBcPlCeviMGP0ZjaJLdClY2p8iFzLHKNmNI1YMx6vXICSfxMSqDqE9/dpNgHO16bT9hus2RhFPNB2
9jfXzkYvQjdciDYiEViYHZzqplVUdgx2GoZRkyBttr2tblYDktFe/t3cAITFL7y/vrJZhUcLRzSciqHyuJCSFAJb7yLsF9xrDCxLUER5vxGBv7nNKFg/pWKVmDU7FcQp
WLg0iE6vTV5jy7AttSxz7Fw8OIgoER46/ZZhaJDZ+Bl7BuI9M77PL+25uZ0Ra7wlGDkhknwdndRBi06iyxGbdyOP+d5R79sHHyuDpqG3C0GDu2Iisbhdn9yp+ULj/dL6
lcgUJpJTsJCtSOYEELbc+pw1d/HYGLiX0yVbwBDnKWINhZId4/NGjayfClB45a4JiLY6/J0doFWSGkuk+oJcux5KlGXRhyec6Hiu0N4FTFZX7D1el4q9XQ3fBItRg4/M
nzhu6yNXfX2z2J4T6eD12sO66AjIhpjHNiWDGatkOHy9nxoIzN553c0QgK8Efd81Jirr6/eXmAMKVANjzhtEgn8VWtXhybXXnBg54trEYvtndq/oWAW5+cp/G1kCxbsv
uBNC5f9HkzbIdn2Yst6+usp8MzZymID8RZcLzQN5g4J1NT2ys2xgOoynJuVlTVW8bY5dVPIMi50kxj8CrCcLXL6yWYVHC0c0nIqh8riQkhQh9FTusFksbamkU4xn5VFs
7RisCKWmxTWIB3z5VlXB8cp8MzZymID8RZcLzQN5g4KVX0FXgqb3I35CCg8ganSGiNvFr6YP25Dy9rm95GK/4sp8MzZymID8RZcLzQN5g4LRZTOrlV5KpNQxzuY1u4Sl
2X1Znon7651Dq7HB9+Ai+5oeilK6igH1Jd588E2cnRKXXOTU2YLXEImnDz5y14gcvrJZhUcLRzSciqHyuJCSFPr2pkaTdqs86oodg3qOu+tLYUM/CVra8f1Ea5Wpy0gl
QBr5hWNCEg3AzvysBkRMKy15jW5vrWiDsV5L44OQwPQ5wTtUBV6ba17IH48hlLk9Xg9nyrTG8LbBfMQqmAbK4mCWyMccRrxoR5nCAHnqouhLRkMEA4wwefRuukZwWJ46
UyYjyPeJ4g+p1c5hoeshQ9RGZhQ+NGo16EUA5SG8zuaTL4HXQ/wlvq0pwe17UIZzJPzwSHOxruXBtdwSxb8bjdtknUGg17jm40blznn8JHzKj8wRHaCbcLxm0CIzvTFo
0Z2xG8tJx3rAu3XcGVDHai24u0N5UGkmqgihDsQZ+XwO7wwTWc8XMG9a9dIp6sIZDAdc3i5yFZrepXZBpbAkV0i40CwSuFUriedF9tZWX5t3SVgOruSKBb705R5K8GPF
T5Yfw/nw9yPCC1tBgs1Wi0B1Vi0pR2gUXSELq+1i4SmhjBlGrU7VIED+HearoOYPFrJzjbPAUTd3hJHlcsbizZ0bvupPSkv/bkE9dD0OoHLFW+2rwx0LrqGauMVmKpty
/ArxS/Z166l2bwIqCG9P+wO/1p+fmqXN2AAk4K4EBxVH9vfPP32vBDIuLogmmGDdFmwNzLH74SDH8apHMa9lx9mMHL0DlafbNCJUaaFG9f7Wdj0vB9+gxE83j6+UP2C5
eJhaI93iYG2Bs9IIVGqasRn8VhRqUKmAvl62EObTRtawmPGI2Bxdp9hmRTpqzsz9K6PMlmDluuVfSOPvWyYFxO0ftegADdiYodD6osGMX9XlKuv2bZ/udZtZkbDBuBzg
wV3kb2eLu7Mg345oj2E9JTDWTaUyAvX+UdtO+yuW/LNf0JA1ypW4RKCIrdTCYr662itrahyL1QMT9kY5ZV7l/tBwjAuQF4OT7pY1JPdE5GJc87IOTcgLSaToZt+lYHjU
5gF+2dtgT7bOTB+WRTtMKMK2lpHSHsG+F2PFCc9tC+5Ng35foalSW+ooXbW0Wj/umX+eIbaBKXuE36ZPKuNdta/9sBT5mjhAt4aE//sV4EB7BuI9M77PL+25uZ0Ra7wl
yUTN/5JciyBjzb4qVnV6O86v8jPhfoyGcMODFknA9RRg0agPvkxw8IHVtbhtRby9l0t0aX/LWzEDyxnWzLGZfRRohEeLkrWPSRsNwhsVCRYiueEr5TMpMFgWZLCIgE1D
c3T96zhdCSScRzzLZnwhQp59DruMZxqVkBfVybaJiJNrjkBAT4K9Fu0Qt/XM+emiD4TZzeWWO2lFEsKzNZtxTVDhScGQMisBMGbux7SOpXy4qXUqP2jj1RpfGvXO1Akc
XUaJAvV4cOYzacAx2tyVnrb1aRqCVh50WBDzhlIeqeVr03PWdkO007tHX7mhMB2NxEpMS36PqDsd4tazzkKwjKBdlqxBZQ+9kyxH9x/V8KxAOycLx40EyzLtRpAk+ct8
Mv7JoGGBygBDFxmZj8G9hCrKN1V4pZnsLk1oKldIysBr03PWdkO007tHX7mhMB2NUtm/o1JJwghf7H3y6zdh7bnQgsk+5onzGLGJirzVHpDgLY5vXwU17u6A8iKMLAU6
EIks5L4eRsP696OBQBRhwfmXOe8MslHPV0pZLl36vyV4QhPWcu5MyZmcX0Z+PNUjLmKRiI2lIu7X97POMWrj6+KDWBXkA4YwMNZ0car2z6BzGvIRyjPE1IuFLdgOkVY2
j2ouzgz4UN54HcG5SeH4GeE5wwveGCjcow5mKkOZwoZzGvIRyjPE1IuFLdgOkVY2j2ouzgz4UN54HcG5SeH4GXY2GoLfXzO8TbI55Qeadln/7ZdDiLWvFbfFKdpVe6lQ
lyUHiuskb/phONJWWbYaZhpPbCpnFJqtEZYbHK7O8t1tSaPK7KmLrwyxNrV0IZnBNR/MzNbjumL21INUdvKPUS0prabbN8zBdagKQBdOqz1PuuVqDwoIGnsrypIctHnS
UCZdkzTQm9xU5ueQUyKGnlSAQNX45UhpOCJd/ar1YucVrBPaqdngUHh9lZuLIhhE/+2XQ4i1rxW3xSnaVXupUHWtzjNivxqli8C80+XJQdEiVoC0ikdE2NhqZrFd4lkj
G50xSk68S+Jf6kO82xsWSZS3Se/7fBzmLnLAhx08H2sdDzvCjNT77i2NpjkAPOm88TJACquivadSPetcg5sAjg4RAFbaBHQjBzhiMpZ+Gw4bMngK3opv/gbuUJCeiTq5
0kxnjm7O3yvR/8xOiJwUOYvzsVukaGa6N1yH+UEpqbUDLTN4M0sCup4Fw2v4iYmXuvCnK7tKLGDYxdvkKcWLAZRobHU9JoRxnqmKJPHA7fIreMsyUcDMG7T6frz2BeQR
+RfxYKXWZQAenfOjKvf+cVoRHqAhd7NP22EUCgf2JAb8zk8AewojIMyBviPrlmveoTyj8ZSbwZhRR3qCv82a4Gn8zpLa/Xzd6QutQ6PdTdhz+bbf8X8v4GpJLCntJ9DO
yogm0Sa9h4GMq195YwJtiI9Kav/JzecpTs+Qw8Hr1/Zb6Wsa8gpw3TGd114w7L7qe+2GCQVTbpRs3GvanR0mNJIAv+pmEUB9yKO8U2J6AAvU5knQzysEZGbdyKjfJ9yK
jsctRrp0CoM+Rygi50UrnZgTfLqRlhv7pRWcHmpXldLYeiksBDkpt91ZTCLEFNcLa6hjw/rMqA0OEsfeojCDpAEfa3nhlLq4a9Hf+oo4IuOz0TJzr3Adi//v0lLzCnZb
vc2DxPnBxd9/9l4VqLAYCD2u5hk0Qpg12dl3+TlBb3WwV3yNnFeC2/R35c0XWImxDqnVP/gAzl+xxt4WrQGd2q2WPl3UpB+JWOqJkkljU1dPto6TLhwOAQKpmBzT0SSd
5EO9KukrlxaHIpWujumltFGi8K+QXQ+b0ucrpT9/ntMMAdsx1HhGNL+qMJq59Vp6iE4e92EocfAi5Od7D8yvPlGi8K+QXQ+b0ucrpT9/ntMMAdsx1HhGNL+qMJq59Vp6
jhhxb3XT2zZId3bdkp64ikTHtIO7IXRLkgBzXAaIVwmslVtjpTdMbwc2Y/VX+Ma6Lc79V/vlmWO6ofuCX4ouHzbAl9Cp1yvZde7upGGex908oQBKZQKIkOvhVGr0FdDz
rZY+XdSkH4lY6omSSWNTVwwB2zHUeEY0v6owmrn1WnqlxfjkL3igc8uQlC2fVkJ0e6KmRNvqZHrEfyXCYGSwmAHtZdDRgsZDWxtVoaixms6DZ63cvbZfXkCwfUipX5LB
N7iDfgqKSBZM9YO80p80fF2ukQl7x3Vn+XUON7GVr3kaSaPqyybUUCnaeNsuPxZPW+lrGvIKcN0xnddeMOy+6u6I7LRzLcd9WPL+WSO/jfcqQdNgtnd4VWBHoVyrxvys
hhV5+aUXWXxZ5AKKr9u5TwDpco8sf0PlSuLNIJr7x7+UgGMwBVn+Ro0ZQCQacSNslZuWpx1fQ4dNYU+9gGDrCtTmSdDPKwRkZt3IqN8n3IoRew1Yc6FTrFQcO21zw2su
SEVuO8AXoqv/9vhVqNg0o248f0rtGQN4J7ofDnxZ2fWShFEPum5NWjpCgqaDqsAB7Tp2hS4dNwQ2GubOqiYZZE6URw86Myjr5TFjAY6GOrQoVHIKMbS+apsVZ6zCe/um
r4OVlbhEWo+bx8U2uXNJZEx0B8eIlJ4kA8PwJ4VT9pJkHu+RYcznWWaGKFINZJctZdrPGbiOzipjtp7CqcpJ7XaLK4uAPjcpDNaQjnEcIyLGQlUxQUms+pUUCLmQDBzh
9K6IqKqjGSf1ArKU57XHP5y1RNKoNlI9a8LMZU/pIUeW56J7Bj/1CNPZqddTaRg+uTHwpjj53V5y/Tsii+KIBTrS1FrUozDZqSFke4wRxfK375WKmbYMAoSA3cFw5wVe
lVvndgWC53OYF6ILazncuayVW2OlN0xvBzZj9Vf4xro8X3KRaJosIafJQ7Z4xDU4WCvg+l2DuPHF8Uw3szYwj8jRkU3bTUQvx0QwRsrrLBQZlOQTiijDUBffYYf8U10z
fLIGkjpJwKmholowANhM5SUQd89Y9OXdpQqBwpfz0uygoN5MQAr7NhsyqKsqvNoRdWFuYcmfms28Epm0aRm6ynFFhFzj6ef2lptKw2GKkJuuV8MfELhelOR1Cp/+KjdA
1nY9LwffoMRPN4+vlD9guQWhApW+Fn2SszipHwjJoa6y/Y56gfsA1gyBP/JV4H0nHV0TkCjiM278+WswTItV3Z+6aSL1iRO2JPTS7nhoahxf9EdBc/IG6/aJYdO58Ca8
UKXH7LPL9UN+n3D8YYtv0apmB/VKu7S+Ay0kh6oSkxvpBZDnOpaTc4WdvrzZe1cMjMGRJzlB5bTr3zm7lFOiqsJjCPQAgdn7xw/zrkQBQ1AE7xUYpFoG/PvTn0kDvlaW
u+aD5l17yzwd6aLpbyiI3ToCAuaRBdmeztOhfULZgOK8KrU5au8kYFEBP5GN92N1Ns+VYRj0vJjm8rcE4ogFBxfyeqgItMgX5EjB2sbBYYNQRcEaQMHC0OG1hScUsleC
W2q6gv0wlxsIoWqa469FXoxNIC68cUokBxjrq7n/flv2Ep5WkTgLnEHmzE0Yd6l7SDdlM+j8YNvoYLZObteNbHZbwn2vylcszwKTC/JVLGQAa3auGF7sdhWylEQ1C1Fd
JmWZEzuEvcUCfO2J8JmAfrWKnzJmXzsd/K9hBHINNBf8TFRTSKiTDQXnNxBQVnvz2aSnM/blF6PqDSZU7BFQv/XyRssO3bxm3tWVTrPlkqK8KrU5au8kYFEBP5GN92N1
Ns+VYRj0vJjm8rcE4ogFB0+2jpMuHA4BAqmYHNPRJJ2kzClCGoXbWtM20TbCxsiAZc4H2GOZ4qx/SfTSBsBxyvNVdTMPLuDTII6axeGqbd/9P0tXiO7nf/OFMQr4uvWf
lsrn6QmPF9kB/qXbvE/4lgHLNo1QvMHFh1eejoXg9Uv4zVZrOdafSAHCdMQzUxS2lWeZMokTJIg6AFoX4HSGaTujkSgGXCXmKLLjuRoO0s/NJ7G5NH/R7cs6Xo5egbQ+
d/rWwK6V1klySnH/0YDWR6YsQ/Velr1ilTCaLbJK0H5BF1oDnCZefgrKjpIoOCnpTZxHWgbxy8Sh+saDvE10NFWQ5bWtSLFNWFlWfSQK904tyL2NSUq/TkgGRy92LEn7
BXx/UQRaD/yXvqUA8Nf3r0g3ZTPo/GDb6GC2Tm7XjWx2W8J9r8pXLM8CkwvyVSxkt1dQdNQmCIMw+eqMSwNW5iu4zXpiZxuRfucU1eOa4fprbgjettr168ip2EkOfGVy
XJPqACXmvxdp9FnIDc5AujifZ06oIe4/xoDvuN+IHt9pX/HDu6gv+/JqhUSDjPZws2A8NcRnPE5xOaV4ESVdbXGysZyrB452Ihwd/JcwgoOWnTJr/9PfS2jsaIIAZ93V
Q+w01OJJfKh1N5LQB6682AeiAMkSsz7zXc2EoMlPd2SkOQM0e8u43c/bte5TKAF5jTaIMNxCWIZVhvSJmLgvTwFzDg06VI63Vqm71YEuQZ8B7WXQ0YLGQ1sbVaGosZrO
62QmMlXpBz74l2f1qR+AeXHbvvNptc9XIAnqCpOornGqZgf1Sru0vgMtJIeqEpMbWaMIICQrjt2koM4qu6YUPjC8/owRb/bFyJAqOm9QG9sOnMNfN8086SKmGzUI4Rtm
KSrkrWY2dCJ/z0PPp0tkwgzBGFNpmgcHMio5iQVDUV+SB4StgB1owWojKsYdwdtV6PIlKHdr7MTk25PtN9BYbcPKev4calqgLWvkl76TchJVk8VtNnZVMjkOEXQJZ1VA
HTnFHdGxhoeWihK7OpIxH2BtNSEPaNwogtvPvySMRDtLFgg4hY/FMy9ai5vPCJ4uJWBrYZcWoEnuz6nPJ7FipnfpOstTIVJfBJA8QZTaa3MJ/2iV5hskkqt7V74zDOv1
Ku3qQQtJi5Tjk/k3i0WpXqm71C9ffb1f55NaPn2FJ2in9lgP2E4K7lhUJiFcuzcBqAiFsBwMgBtoaRm3YtERU+7qQoCImNLRx2gozVdrxEuio43+PoE23VgfyDzcmRj4
Cf9oleYbJJKre1e+Mwzr9SRaXWhPyIMWK2nDY2HcaihEc0XXMWug3BlI+MnkMqhmOJ9nTqgh7j/GgO+434ge32lf8cO7qC/78mqFRIOM9nC+AeuYDBQdPrW+MhAcqvWV
POu8QeemDNNBELFb2fPQyMysPdWXIXfbnMTuZkxcRx2F6hsw2B/QqZFAAWdSPdcnXgf0fdJqdEvM8wz28j3c1o+oCLiY4TEtcZuZprseG2WfW2q8nEkWvdp00yS3DAUm
p2DJlG7YNkbFH7fDbFz2bQ04ClfpDRdAfoD4aYLYc7lEzUHyiaYl+N1T3/g1/OegbBJcD+9xqGZ9oKq38M6Oo2azwiCXU+Dfyd+14zhUUtXsn3XDVKZN/PkjvHetaxyW
UAqebedyrJGSgQSkrHLm3zlDtb7tZNitdA9h6fESB2E+p+8cqRKw3XD3WtZQkru03osZCR/Itkbv//FQO3gjP7NiUP3WbggTd4K+avL9zVF5sPN4FbyQGRZnxRbDt1iv
i4ErRzEdRuI8GlPc9TwOeV40cql246kSm2sz01pnaD2zYlD91m4IE3eCvmry/c1RZHgKd+3gNjeeP5glZRtRdYO//OIC7ed6nYWhv6QNLPz4ifEzJznlx3Z2WQb7cxm8
r3ZaB0HAX9luWabs0wTo0l1UKmI6/oMPxF5O1qiLi+mgXDB4s8pKeEkqh1JV/Ca7VAGlGb/Ybrn9x+ex6qdZTm6F1G3GU89zWtNwIiPlnRgC40AB7HnSUS+8bclnkqO9
EvAmQbsgaj0Y+4Cheh6GujUkW76Z07NMOdBg9AtabKObpZZ6r5N6f6QKARIef+w97v+DO0MQPaFaUQ52HZ79BGlbVGW3kJoRUDHcLOjvc10ck8AG1N7AqPf88Fn46msh
Ce8JYDxTXzfUrS4F8fAjeu84jN0i47sp/JJIU8aKkDr9lQMvihlcA2gqxa4WcZjLa612c3q6jvYKepM2p6PEdysLO2XvjBvCu80b5AG8/VXBJ2EHuOQA+iFeb8SDc4Qg
K7jNemJnG5F+5xTV45rh+sqTaGNjSo2QfiAeHt97FgXemcgGPr2tRGVyaYAroofu/aOLKgDCRi4PPNw26JB3VcGNP6bVjQIWMDKg5P5j/gkLR3BhRgCy9hN7F+yQ3fhO
DHV84qRdlXAndTLNU0AvxspmdYEDs/QOxx7/ur2Mey//9wTZIioj/h+sXupzUCd7JnkAwbXSzCOCcH6FOoiJn7NiUP3WbggTd4K+avL9zVHU+WpY/XiKi93eie2vJx7i
UbsHtvWJJryrZbpwF4rWcSl3n1NJ1oqWhhhq9hsA8l3ZRFFvd7/RTibIx3assUXIPm+uhYIBIqruXCZCdPpLbBPxYDyeQhfaIXqmCkci3cJPto6TLhwOAQKpmBzT0SSd
k34YB/34yylx3ToKuvEP74ZuTzGCY2HKoo9P3gXO6MLcDOjmtYCGctQcQ3ljm44dXose9QGBEsLYCcguvshtQSmmb2teqwEAQ0qdFCJvyWsxpRIw7V6t34uA6/E9M0ud
neuhzoQKyWgixSiK+9gMLFBBtUcDFefktYlvaa9owacGnqf9a8oXQ8r0iBr33n6bT7aOky4cDgECqZgc09Eknd0f4V6+2kr6Rf3t7YDerh2Tm8Z+k9iPQ7CrUkGrBLq8
iZJhylUCX0xT670zFH+AvtwM6Oa1gIZy1BxDeWObjh2rnu+8hunNmqskU48U+l9hmtJu2HX5tPEIsboy000TNj28T17OhszgRVPJ6Afu2xi+AeuYDBQdPrW+MhAcqvWV
+MKWs9PIS9Vg4bYPQ5yvjcYW/aT8wSTF4wz1Lx8/j/eYRhHLkcc6X9+/qmVBLFTzkccEjCstMd6hKeiSCe8XTQ1kcUe7PMucfvvT9oiclX5jeks8acwQePyprNkANh3y
8U4HgspUwBAw/ulm4a41hx31I2A0ogt4O7MhND7oXUR6tox6npPn6JB41lj0ozK7uS9wqOx9T0hST+VxxdddX2uEnJTTl3gVs7guh9Wl5gU1l7DqDSHzv+s0eQDC2EJt
JJkPyJxyLJT5Kp5mqL+ri8y13KeJwLIbOoWXS6NmoT0X6Ml7+BZS4N7c41qTW+jSdEJlt7h1J0NCNqOOWJQV7oCAS7L9YrfhMLpRRCJyRcOL7YWaEMaV2/yIIywTto7K
+J9h+KovGBMCYQa/Mj5O91XfoveqvLC6z1pt0Ijg6s4a4GA5CQIF7eHEJZNf2pVtINCra0ICeLYWqYC8KRGd3jnIkRvUnbrTzjzSU087DvLS39wPAxTAkKHH5V/BN+gf
FrqkgyE0thwEU7ljKuYFIxpGt9n9G9foTVVrfoWs1EgJ5Nr/AyuveAi0t+0V2Cuebh1mQOz9jUlnNjxkAqdICDs+FcowHIPWZY/nMBcBQ16N34yCw4W3o2k+f0kSsKGu
uASV0O9EFGtPqbhf0uJYJWE7CcNaA4U/EBS9KodgHwGB91dGaGGjdVQrgck0Qqx1HQ87wozU++4tjaY5ADzpvCJ3iJV2xdZTZAcKWlfEU1pShUVwpV8PFCAjDXXO//+G
DYXO2Q2q0tzkazFEYcun6JvYE2HnlNCT5vyDAgXs0Wm22Hzp/bvx5xqd6ytWejcZR+sTsUrmMdAwE2nYERNotoAVFwoUFuI5PVf+NIlC2I0Cmg0K93XTTXfq8MItP6eH
T4o+ycFjNLai+e5fFZWDz1UGiXUi6PolPRZGKWx9WFeShFEPum5NWjpCgqaDqsABcCfJFAXFAN1RoLhnjzfRSCTSvKz+W+VPf6U3Py1Tn2woVHIKMbS+apsVZ6zCe/um
WuEiOdHZkRf3lW1reBJnzAjNjxZSbDLkWIYr2E/C8jgl0T5RNnjNvhZEwIitSVEd9Ou451R5mm6yUZqGcAPCZrmOc/1Ih1KsLB75jq5XqUQxzzZNYr/n4Aw66sYajX5L
zAfvXGnYjp5E0NJU6HLxeqx3+WamZUcDxJhYUpP+wINNpUKrSowCUN/SE4//3wvPONjSm6W2Jf7AQ4IgufSzJTbV513lc3/eEEYp5LP+NBEYKOQBy0DE8oUGiWWsy0fD
mefxZdZYDa4W/IZU00DXKH8+r3yFVO8kvZ6qvga6U9v2fq7q5J+jzFpse+obl2JynlzQW3r11+RaB+HzLkTUDC8jaZE2wNcsap6bFWYEZ+oqQdNgtnd4VWBHoVyrxvys
KkeQd3JXxlheOFA4vMMYtkZ3tboJX+q+FgOGrPhjdsGQ3U9q3FAufoBEPwYYR/v1GCjkActAxPKFBollrMtHw1omm4oS288ZbdgbkngcbgCuyCcH3NKNi54OjWYgXTg5
W6AMpoQBQz7qlyfBccrzCuo5Vi2b8fsC7nXPV/7tRhAD4d0ba7Dmm5fcW9QMWGe6NknE1sRqzoga8z1K/Y5Yy9VsgWI9abNtiiBxb5S5xe/0B7aqoIsuzQu1WNxDcecc
dlAqspHIFv1SfrEmtHTBpno2Nt6nbBDhhtYlqskW5pUFcetbs6j8neFFPqydZH007MsXxfhOvGwCwd7b7qFVkkZ3tboJX+q+FgOGrPhjdsGQ3U9q3FAufoBEPwYYR/v1
TFdy1kXr8gcFoO67/R7q45hE6qMC298qG2772PLtIiIt3w96vD9gxah+rxUcccuaD2VaiJf297bN4fo/+0GDvijel7r3Yxh4yolo7tAs6tZdArsb4qqR4InIZbtqhZ5e
3tg36JZIjTN8D7VQ9R/VspMJKcofYI88ZXIKeV6eAFkiuhgNbLQAA+OYU29OhpRGKkHTYLZ3eFVgR6Fcq8b8rE3WEGchrfNfvj7TXDSATQ5HbE8R0jHvFGkRAPbPyPGB
46D5UnZvjRRFTBDE5JM3wETHtIO7IXRLkgBzXAaIVwk/CQnWE7Dip3rSjOnIwjCpyYvCmEqDqPwxC/GJ1CkhezSkrmHpfvGKFQ47udGA3Mhr9XQ2gbxmXL4skz/UMPEG
6CUPxBjAyqLWKj9tQ8RTtysqaaYwSOA9GE3Gy4OmIdbNrhPxolzl0CyygTfP2TzdjM5+QAcLFc3Vc83HAF6nB9Hd3c270GqDpL6VWmdXKEKITh73YShx8CLk53sPzK8+
PtnXRYZprKsvEaCeB23x+rBiwcIShUPnvDmqngomVKniZM8QCeDDMV5PHeVrbyLc5vkjfWgnBhKOYatM2lRr/kUbocS1NYeMXz4geDDdQxxCjFd+OmdLCrTQNI/q7Loe
B8lRZBoeBsWZiTO6bLjcMs0VXA/QfsMuB7uceA/b6GhR1K6352JQ5BqnOT0FE6XD/3vQwyp8Mit6vANbO1OFpudZzmN+OjXTp319s/6X1qv4lIqPTYIqr5rLAVLXc5Wv
AHJgYnetRbFIpFaSqRNcGjDNOswLA9rSdRp+HZAEsDZqSC/tqfsSmr9NJ2et5TaAJOnDtzmx4P9ep7vNCFhsz9ynGNtO0SyBEE/lnZbnnwL6TKnsRDdUgZETqEJiDdrM
laVSsdyJi16WXcKZbNgidwh8QdlZyd3MKp8oYsf8gCAAa3auGF7sdhWylEQ1C1FdJmWZEzuEvcUCfO2J8JmAfqJmFAMbWO4EpX1RzXo4TAgijg/poXCHMImAxGusyuXM
pDkDNHvLuN3P27XuUygBebF4HVpgESGnMVkF41EsMcmOC88ABZf9UzRlnaUbdHUXAfgfD+XmAgw7rWKZZemVToGlui2WFexKAXaUEnl4QXSX0+goEAECl67ggp3rXc6T
a4SclNOXeBWzuC6H1aXmBZ6Ksz8BwnJ0Dk47GAIwWh3o8iUod2vsxOTbk+030FhtQAHEcuUxEoqodDyQB5O4rU4tlS+3fA0QJpJdIs/lM2yRt8GppsHjPP7FBIuQH+wX
pKNR1nfsfzaKv+tGh8EOthUhBb365eBlIAcPi8sxeaXpsxCkSiu8zfBo2Xi/lxiG8pVBoGJ9QV4hfcYucX7uDFWQ5bWtSLFNWFlWfSQK907AvadNpX6ZoI75PcZlXGBk
salIvu8wbo0t3GAwcIpwTDDNOswLA9rSdRp+HZAEsDY6qbiZxnFbs4lmTlVrExIh9w3/SRMZ2s/eQqI5AaxamgOMYQa+ZYIYSbu/jSFAVhqrSpVVndq0wwXXZeJSGUYQ
swpwncFlSK5WfIALZDnftSp4sQDDxKAqO9Ik9WKtYeWgJVS5OOZiyS4t252Te02fvCq1OWrvJGBRAT+RjfdjdTbPlWEY9LyY5vK3BOKIBQfrNLH/8eL0dzgWkcGkDUve
41ZhZuiDJiyQK2gC5Qy4p0fn3Ag4CkFdEebblBZocvnZT5TP7h+9AvtVGqrekbPD62QmMlXpBz74l2f1qR+AeXHbvvNptc9XIAnqCpOornGqZgf1Sru0vgMtJIeqEpMb
gPu50q+YuuB+Btsnfl3MPgZ8fCjQeQINiGnuGHYu1WRrKCqfk9nOMiVA7n2cM84g0mjw7/vTlyxhChotZcL+YExXctZF6/IHBaDuu/0e6uPqVGxhX1Kv071PtsgIVBlu
zKw91Zchd9ucxO5mTFxHHZHeMDJcymm8/A8ywtb0b3gL/kBxv+3+pSyAujnhYZ5BQ6GmgBQejmTfaCJ6Saw+5kvAmwf+gE1Kr9WWwl7hpxyDZ63cvbZfXkCwfUipX5LB
sGUr6whSXs7Fnfq1ProSpVWQ5bWtSLFNWFlWfSQK9055TCe09TSHMDFh4f1JrkDihd6rsX/CEBEaA3WXHNort9Z0iGkN1C7zKjly8+pHaw2io43+PoE23VgfyDzcmRj4
Ua8e+mBdBZ9kP+oa0sPh/uHNPTvTyNgd2xn+yQ7LFS+UUvEQlBpyde/UQpRwaY6UUnUA3y6KEywOdoaDLiqkoVjLaFY+l3V7vdkikfEJUvZrrDf+MhB6gC1M42QI3Tck
8p+GSi82wH5TUsx43dW8I0/fDQ//nh+2JwkrjZSLmYjr/b5wQL4n2DQXTuL+WJvjWCvg+l2DuPHF8Uw3szYwjw4XUBt0nryBxU8YU/aVkVDbpV64fytt18JkuH+U8Lwe
DunweL5KrkIVNRw/yA2mKD7yt/XGYOX4nhrLdSBZ1g9j9KxNaWYIh9sSYDxy/ihMf/yyJUJ1gMdgDKizi2y/5rYqfTTrUDGb3lZKrtHJiGTchhFDbOb/09bE89ETHk3q
FDh34bnR9pKxvkwjOdDzq7A+rKIcOgoiPEBPYqcAkg+dgh87pR4YqJD4XY+De5BlsveDyZQfdQarv8jHEdWtrT6wkhFUJ6SUVlVlsCY8TK2G3SE821jEj2s5QOq/U3E0
SDdlM+j8YNvoYLZObteNbIK9Cc2pBoqSEIzeInLeeiM8IvEL1AeeMK6HP91TCCFXgJ1gmOBwUWkujoXPkVT5AO2QLVmwnlRCOsgqroFz9808IvEL1AeeMK6HP91TCCFX
z/SIuci6pm2CRqDd9nedFW0hFbXn6EgJFXWi52UO9eaqZgf1Sru0vgMtJIeqEpMbF5t+2aGm7bPkXIGIt/U+B2gV+pBeqDBZW4k+FCS3FZ3AsxWR1qYpty6iQ1ROz4ND
r1AZ7Ta9eOPTGdMu6UfW5jKVI40OtFdp15GOTDduO5HOsKGRaOyohvw4wzVTySYcAsMhhyAYzcGn4rTt8cBn22AB+NTV/w1FlulJ0nfgshQ8FooWBNyzwG9uL2vfz/ay
sd7Hgno5BlO7Q1dP6rwAMWBqndvZfAKzjPxP1FVgsMfToXczIOBi9SNG+sRRd6oQFmQLs0t4wanGCzqCMf9I+1upA7vvugTdGqrZJjoomv8jDD42uFVKwxUUWJ1+Iyen
RFnwlLzKCVGO6IONvqsNQTKGVpAS5u4SzPYEcIWxB8PDnzXbEnhyM7GIeSfXUqyYqL8yhZjeNPODdF5jTxxiNMM4BQ+JACkMlSumf1qefZReeKOFW4RcJ29CK9vUC8Uu
rYRG3pe56FIdAIZvmqBr0S44nula2BL8d41Xpp1gQbXzIDqgy0iU+PAcNZH3SqfAMm+ghCr5ZMIP2X0/qj/dhpTRLewf827hiQoLB0WsZGaaldS9bTTK3f7HX96zq4Vd
LyNpkTbA1yxqnpsVZgRn6rS+gEIREsHOlKS+DIXPV7DOZ9PnTyoql5Kl3m7J2mrT8r7SOloffPp/pv9m0MAN1fQHtqqgiy7NC7VY3ENx5xxl22r5jAIjap2RXUQsaA4I
TSWS3j2NWtoVD3djky7mwuEVeYBtHot7eYFbO3lBiAGZ1B8rYsmc2DRIWT6PLmgSBA6piTaJP/UcrcWZGse9NbPqzge+g22Bp+dJaQJvBsDtRDWRUHw2b1glgP0LxM0D
2/bKtlshAIdjfLyduhFtRmfWk5t7SYxhWWKXGkdew+55ess4VS5XF7cYqIZAdIfzY1C6BWVRtqYcrvkWZ/aqXFHulD3NWwXTpKWIZQQTPoyFWNRKFORHXfAtX85UQHs/
WorFZiZ2n3xSQOOaTQ1IEM4oMBFFDYYdjC+GuuT1X7bCXlapOVkTDphEyAOb4sOU2RSRGFSm7XHFhiZdlmAk7SGj9fhlRzS3MEzRwWlAjtl0m4EEG9mVJ17dWE5OAOZ/
JjJ2lGNEdO8b4WOU1p38sRS2moPKznFiajZW6w568TQvU2vGNxGtBfN0d/sPHqOEsZfC8Dfzp65sMj9kzJj2U2uOQEBPgr0W7RC39cz56aLeMM6nToeUKbH43yq37N+M
KbVwFv7lmIE483NxjEeS0YHP9pyCIsCdfrhFFdhKxsQApGqra4vtO/o+ChHTWRwTVdzY3EiwwpZ9Sopd9kQ/pKh0g37yqFPKzXnBFVLCrSyYGD+uzpFhfEYO+47pMmvS
1cgtwNMgvuQRs/yhfkjB8KjOmPPoRIN90TzPv2pqPoDYcRi7Bg9qI+gdnegW86j1pXKHsJV0YqrkbXM/od8iOhYvw4vThXv2wHfM6DxSWlX1moZGNTlf/ZuDuRsSz1EI
AmXIMM7kU43rxJF570uAWbDWg+vmv+GG9zVt5X8FznArdD0UjviTO8umh0gr96Ylysd9gvob+ltQc5P9gpD7HKMUCeakOP2AO/yQrYJ0euNvZz8WHCAWbvpxrKsuEkA/
qKMyKVtAkWNwlCx/bPsBK0ogazM7L0oI5486ec+sUNEI4xUcBOBgDvurw9Is28JiSHU+DzHHUlNkOSMK6EwXZKuxgTB9nSN4nJkv2XtvHpN4pemrj++X5hp0Eon7BHgj
jNrpVyXsPHTagFxhxNickZibu86hXTqLw2OKlXVQJjgumVv2Y3sTCrkrlfRpe9eW+J9h+KovGBMCYQa/Mj5O9741TCnbi48OkR1wMCbfo/aTTd9zo9gXac2imlfVhkL9
uXru5oAvUe3zoQR6AztI8loQcsPzgoIRTmyXQQtfyrVkjb7owkbC60XvVJHOWzyUlE69KjbZt/kTLJTYoDAkeU3rOJQRgr35kOQFvB3frU8EN+MZn27N8v9Vl5flb4h2
YXnMxmV1zaAAS6Ugesp4p2SNvujCRsLrRe9Ukc5bPJSpdDfjbTRVOdB0wgB1fIXaU5sfrIsuBQu+vYP36m19UAQ34xmfbs3y/1WXl+VviHagK9acz1PID92tyXGCqgmc
1eLC6Jvhtty7WJfRMxP+ZNQ0YVoNsU7aUaS9/300vkrZ6fo9rCU55BGXqN+boeUQ62OBnenKG4C9JOvIDYwNau6wrVkxhOLkC6DF1IAhBbPLTQKawyhWTq0qzQZ12mUb
8IzAWE7NTXEEVp/8ztQeHRCJLOS+HkbD+vejgUAUYcFikIekOFqKlykC6JHM13jgmFnp0MCX1o0ZDe4MQ5wpxTkJ/s9u7Gk7H+f7wRicrMa90fb/oxMiZl5VQK2USdYo
WAX0aSq8jdPnfYofg3WoHW/LcS6c6qui1mJ57qXDDaCBJxHb6Awuf8IUNhAWOM+a47Ue90Y+g/h0xgK0gLZL47bLy+0QkjS11KbpKhvLCQWb2BNh55TQk+b8gwIF7NFp
Tiq85gLni2Z3Np6TIm9c5FBjqhObQrj76C14nS6j6XodDzvCjNT77i2NpjkAPOm8n0ffZs9+wWBCwzI0Nz6khTs+FcowHIPWZY/nMBcBQ159GUpigm76lzXgMOgOgpjU
WAX0aSq8jdPnfYofg3WoHfmQDAW0Pcc0Bzgy3ea0c+ZgITTTfUJyXk3Y8vn4x4/9kN1PatxQLn6ARD8GGEf79WwC81YJkUqczhWYrElGThvCeGlVO/DCgmv9+0YTEOIT
9IbHN1Yj7B5WhBRJ9PDbvswH71xp2I6eRNDSVOhy8XoIlhi16nOyUbFjGju9qe/CHmcEzAtP6wSVwuUCrOrzcKCSOXXxiFgZaWoV5lpWQRC/fIivdmxzTEamHAr5xpJV
KkHTYLZ3eFVgR6Fcq8b8rESyf19H1QH64eVK4Xmg/i5HbE8R0jHvFGkRAPbPyPGBFyaysOzC3qANVZAisEYLkMqIJtEmvYeBjKtfeWMCbYisl9xqJRiJtDVuttUqO7pe
koRRD7puTVo6QoKmg6rAAXnBDymrgNjWH6zLrmbUaLHfk756Qe5Jc4ynP4Fj9sEcQxvBWLbE6DcPmWR9oJFq3MiLbaORSyFYBha2S+2W/RALLFLaTFxY73WsApJEEiuF
3DPKNlnYAsepBfof8W6OP8qIJtEmvYeBjKtfeWMCbYiD4bBaC5hpKpTdxnsQ+oJx49ikr2KDHmwGGOooje69z8EWlUFK0GsQIw5qw1mn6jzN2zbtICS7LPpyY3GIS8JX
n1vOAdXqOVLSf8vedyQWfDsi1kRZ1b9gYIyFla+bVeOQ3U9q3FAufoBEPwYYR/v10rH6ZV4qKAElh9cEJjLX0cJ4aVU78MKCa/37RhMQ4hOTFeWoi3LOQEoviKdH9894
boxlpnbZer/buDSZn4ukbDsorLtev2l5HU3b9YXE7lLagnAn54NtcLLArsZhghW5chamQ4wAWklT7USDJLKoinbp9eomSOgk+L1e2UFEyfsqQdNgtnd4VWBHoVyrxvys
05mtONNeOOP4I8BT1w8W7CJlP4xWqaN0CdZ90abXqBpFvQN2Qb2DvXwanGwT76LVOqLIXIfs1VmZkdhQNy3u9m83ctCJxYoSrRh4A6g99by1l0G3J+2IKlNEOCRgBmWD
dCNfjl7ywjaRjlOWteRBefwn/vbMHuHt/jqMNnW9ddcuAp8gBE08H+0SKLhHaGaSVbcC6Tn8V24xFIMZ8VT/GS5t+XCQVidZkY6XmAAQ7P5/pyfyzQZRZbsAlPU7Syou
yogm0Sa9h4GMq195YwJtiCa8qayw7H1r43fSDmjLEaiollDfX87QrJWnxf2lm6rPnhaGRGK1mP4No8WgMKzZMcqIJtEmvYeBjKtfeWMCbYgmvKmssOx9a+N30g5oyxGo
qJZQ31/O0KyVp8X9pZuqz8u21JTY2QF7PRKRGmTDTWF4IVLUX0E5WigSBL/TF2EYOkLmgbnNAjfIdeLHLaOrhUzUbPbGUEPCWklwWt2q+DEU38T3nFzhbdZkKkt1J4rt
t1p0CWaZhrfk/DR5adN2CPwrSEogk9cq12Fepv4DC6upYh59ImcWLmj8tZMbSOx81opr7rBw28jEONfnWSRomla4FFQ3mJTk605qdqBRjgonCWT4Wq73dx1cIpMAacbI
jea1Y+Qtjxi2t4Fx4ZWdBpDdT2rcUC5+gEQ/BhhH+/Vg52PIM5QL6qHD5K+cx7QfG6x3IFAeuJQ+G7/ycvFRWIGKXU6Kwui6XPYvhz0oQS8310QJ6vsnjQfBSqzqmoyv
HLtPYGZWYjzNDVZIQEy8ZbWXQbcn7YgqU0Q4JGAGZYOQSe7d11s+v8snfqv5EuK6xvbRFVL3Zsn2CxcQTilwHRy7T2BmVmI8zQ1WSEBMvGW1l0G3J+2IKlNEOCRgBmWD
N5BvLaL3G6aqLOT4sjiqBdzXYja659gFM7iImgobkcDKiCbRJr2HgYyrX3ljAm2IJryprLDsfWvjd9IOaMsRqJ45nbXifb/WIl5fHciARJzDdjvsl89VfuWjI7Us/8c5
wvo/qHkmQauBaKco83YGRS4CnyAETTwf7RIouEdoZpJVtwLpOfxXbjEUgxnxVP8ZUzdg56zY5YI85hSFVPcY0SpB02C2d3hVYEehXKvG/KzTma0401444/gjwFPXDxbs
ImU/jFapo3QJ1n3RpteoGhXVKUoHXBysk76tjVY1A3omqSS3waO27TF+le851mCYrGJoAtf65lHdxrKG/um9myoJahreeiCPDLnbr1CpZqdcEfodV4RK7XXJVoq7ieq4
K9tQrzkqtBbnCf3ie2y2Ta2WPl3UpB+JWOqJkkljU1dWG7mfgYGWd3nuKw1OUxy305hJWeQeE+bJZeSbcwpaM8BCxI4pQu+Utgm/5t2LTMe2DqKFDrLPhPjQKbaIZPBL
NXHZLiu+/k1w6ZZ7QcLWDfwMuDL+1UMZBfGCx3om0FZMTYt06ajacT3viInIiXuSLfV0R7RYteOZ+qHf2jv87SoJahreeiCPDLnbr1CpZqfYbc1Gq/4XeK+5AoxRNm3C
R2xPEdIx7xRpEQD2z8jxgRfF2aNa0B9ubYHfjT7tDmZeFFlkoRVezsDC6mQYDdm39t6yG1xsk70ZqxyyGERI72Rvlis0eRrs/OaV5SD7ystTMNnRPzHAdEiviZtwy0BY
GdIhsYWeOnv2QowFnK/KCHghUtRfQTlaKBIEv9MXYRjxSfBLLLfD/N6E7hOvjvRzSIL6MeQs9xMiWoFdMDcOHqKUiIALyV48nDLVES7GDhZ9uJqfGdr3GKQ1s91unS9i
kN1PatxQLn6ARD8GGEf79TGKar66mO5F92y6M4r3c2UwjftLCFbhWKTYtrsKc48NphOSDvg52dDMjZqwHtb4l/hGb1ANrvK4+GgbM6stj5Te2DfolkiNM3wPtVD1H9Wy
lw3tW4cKRNFhyNa89ua2s66kDyDGR0KniNSQrnUOBWIMLP9Xge3hPzvXH8CNGm4E85SnGTRwNVD7S6Rcq4DvPYaX+ouMW5S6HXUD/00h4bJJpUicEQEnuaU4JGmgol49
CyxS2kxcWO91rAKSRBIrhX10UrC3PoY+guUUBut842J3EkF6bXf/Q1hQ/3NbSvciUZ8q+yz32SQAWUEBzAqfBvOUpxk0cDVQ+0ukXKuA7z2Gl/qLjFuUuh11A/9NIeGy
rysRfMC74LO873kYZ4OvZMSgAERSJEJrvqCC2J9EJ+Nkb5YrNHka7PzmleUg+8rLhMQJFAFqoavuYdsL59QRARIfZvIgyPiKMHwBeS0xBYZHwLl1j+Zj2Vu8I4Maq7nC
bBAKYYZoMuVDposw4NVYQ31bMDQ1n+Z9j2VrPCANmKJgXxlb+9c49+2ZE/Im16ZzLIx90vuBySy52uaa72vjQGRvlis0eRrs/OaV5SD7ysuExAkUAWqhq+5h2wvn1BEB
dYbJrNBFqvckdpoJpim0ZK2WPl3UpB+JWOqJkkljU1c5rgVRMkuQJ4UV5axzFHOY7nArRZFQYAdNk1qA7zW/9E8MDui5v3xtWO+Ab7T6cw+3x1tA77ORJz0JMJAalLXL
lzb/5QSFANiJPFqpe4QvOpDdT2rcUC5+gEQ/BhhH+/Uximq+upjuRfdsujOK93Nlun46cpn2PNsnmX9/MHF3lK2WPl3UpB+JWOqJkkljU1c5rgVRMkuQJ4UV5axzFHOY
elsUeewlJvPsZ6XkRllTI8qG60/noq2x6qwFAg8xJXNoY9EPHP3TP8Dzyshya/i6mhu7QjzokDd29jimZE2BylEN0XFVS7qPH/APwydBTrG9YCtFSxohBPK3ocfXLWba
KlutGEbN/eRkYLdZeUFjprr/d6zTt+cL7zyOVXqI7NBN31NwfuplLS5k18eIh3MZX9fk4DzRQJcpx7B5ZQOj3zIkkZZc9dhY/ELIsxkr5+hcAuUM01lxVo/JvmldvAKy
f9Ck8bwkhWsRDco0C/D4QoCHuQCdzWveRNOIN3GTeE1cAuUM01lxVo/JvmldvAKyPFVS5qefGUCjDRjqZ5IvdM3bNu0gJLss+nJjcYhLwlc+cf27bVeNdX5TmCFEk3bk
oedtQEtXEpkOEK5VIKXD1ZDdT2rcUC5+gEQ/BhhH+/UlLd6qRW6DzGV8vnJTgcOSwnhpVTvwwoJr/ftGExDiE0N7gpatpvqKesVsuhtX4SLMB+9cadiOnkTQ0lTocvF6
Y5qKvey0LLJuFK23r1yl5B5nBMwLT+sElcLlAqzq83CpOq6BwZ0xhtzZ4h6QSO50BLfXveJr7OyTRvSJmEaXxipB02C2d3hVYEehXKvG/KzUymTHAtmLWJ1PJoBDMB0T
R2xPEdIx7xRpEQD2z8jxgfT4gbyQmnw2smb/x3MmMzPKiCbRJr2HgYyrX3ljAm2IsngZ8q5EMf9NmM7a1JQqbpKEUQ+6bk1aOkKCpoOqwAHkb9bXc292+GoyanKCYQ+p
XCYFHMVHPisvul3bBdgqPk0CfvgamVFeeL9aDnfzJYxHcMjrEXPUz1PaGzNMqYOQrZY+XdSkH4lY6omSSWNTV4kI7c5nB/vSZUPIH2F0tG/e2DfolkiNM3wPtVD1H9Wy
2C5kFijdYfvTcwC/rCy18uPYpK9igx5sBhjqKI3uvc/DEv3gI7ZTRMF70S13L9SiBbs5D3cYKnEqxgH48+ey2xEDrN9hE/ngfKxo9d7hCLTI74K3rqUldtylr5L95vIZ
3rdgMwHcs5xHKxXHDvdw0IU9iZBGehXFWHStXmXmlA7CeGlVO/DCgmv9+0YTEOITg1SAJ8ctTCoNfIxylg88zcwH71xp2I6eRNDSVOhy8XoV3PPU1q2+xGQHIU92eGj8
HmcEzAtP6wSVwuUCrOrzcPdOfJxHC7v2DM50ug56L7MUDpLbjvxiwXY9Rz/OsUlqKkHTYLZ3eFVgR6Fcq8b8rMIcElbhC0QXr892QL1RffxHbE8R0jHvFGkRAPbPyPGB
IPHBYxq0nD9Sew5mm2aj2cqIJtEmvYeBjKtfeWMCbYiD09fBTK/hO/ieGhfnYrIKkoRRD7puTVo6QoKmg6rAAT6NKyTZyr331yVka6vIAleDW2o3iPJO6jjpYWcta94m
AAaAW32OPyoVCOdwwb4mI2h2obNb+NQnieS7O5Cxd2HdM30hb5jEKszeFKSi7H9Z7pOpskk3EixVYPjUzODjZt7YN+iWSI0zfA+1UPUf1bJM8Jos9Q7DFVI+NnJAQBZB
49ikr2KDHmwGGOooje69z3cXPQ8w3OqUiJkUpLEGeOaHVrkR+RY+S5GVSVoUp5AQLenDhEB/fu2RFLzUFlCQe4NAmKdc6widFnaDTff8WqiQ3U9q3FAufoBEPwYYR/v1
w7RfbZP/mh5J51d9iQb11yt4yzJRwMwbtPp+vPYF5BE3DYKRDkDwavg/pDkqFsluL+QQZSoS/BYqTFTMzbEqF79ZcGzt7ZmPoB2zms1IKGEeZwTMC0/rBJXC5QKs6vNw
ya7BWVj5FyX8Zpx1rPSb1yX/xfdUOA5+LDfDYZfIDfhmnFcOeufM8srPzbgsUi+24oTe81KQyUtCkxF3J4hxU9mZDGUWpO9SSfQdGqobfYBrlM3rf952Rg9E095ep/JX
4kqj8TpC+6NS2a5DiyzsGwJES0XADYWCmNF4JLkeTP95cg/K8OWYlFHE4ghu+rJlMDdo2ohozz2DqCwszV4melP1StA4kYGozSuQnIPSeWvwumHgMilYlHWOB2xyF4VV
h1TjnC5L/ObHpaWuSzv3HeZkJWlyESU8X5eGuYGuq1H2WLb1h1lIIWU66VMqUPdyMHJiHiPYmhhIRa/O9x1SdOccNoybHSFPYwFbwBPclFwZfj5qNGglcvxkE4p352D1
mVlYoJRme2xFmlvyWgB8vr1sKKi4Hilxk6qgeTpVwjArAjjG8nxm8FeiTeAnDVHS92vdDF5C/pj/KxgPUvrSDZJ1XxYpJ4CBzJILILhMHseOLOzNMghKDKne8xZMRxdD
T4o+ycFjNLai+e5fFZWDz8OxcNRmiatWztEYOlJcpN7BrwZZAbTiws17NmKj98u+MBd5ZPuh2Rj3pTsVca59lPXIkaNgSvgGkT3NvAYFid8S/s9kJfpUp7kt6+d3F+8n
GN+eY1dGlBhKudDveJrjpzFiZ/1N++J5mriLX7iVoF481SNbvRUKKYl1gA+dFGT/DT2KOrsT9gjx9wo9umnRP+uQi0Tngin2wgRkzi5Kz+WLkil0UJwP4VVNvOw1v37Z
wgtNIai3AEiK+gjQaW9MeCoMCFB+ono46v6efV+6Zf0try5TkZhEX6fvXQ1a5du7cAEywy5EIuW19LdEMzNZPMy4xvqmp16HUuMVeqjIoI8YNdmbek+X3cKrQEEHH7d1
uY5z/UiHUqwsHvmOrlepRPWjbG+JIKnHypuQ3c5NorbSTGeObs7fK9H/zE6InBQ5EHCaLjvNKx3BBO7bYqcUsQjNjxZSbDLkWIYr2E/C8jgGJq70OFWSlJlM5AnohPXx
1OGiHsldQqwFVKKh01Q/uCu4Jw+ofTu/XSiydpb0YqpqTX3R66rNY0z2YuaoIzHjknVfFikngIHMkgsguEwex9xihNn9f7liy0AUwVcOd29Pij7JwWM0tqL57l8VlYPP
BZAl2k8EBGtOxKqxroFSqQpA1jCWKOunDURWTuzXvRhwHJU4UBrwARIOroK0WcCgPFCiCsciB10GTP/U34fwPR5FB5RUjXttmBAypFld+7w3Z8JQiSiNCo6r9POxnk8w
0i18GYgUAUg3CWCExQYqFr5+E1bl51E2Xc2jWUsqynaTKM1u+2Wg4xOxaWGRQL5Km29O4TPI/ZoVYvTbLC6woJrJhEWKMm4jrLrT624Y7z3H0BhlspJErHatdx+SA2iI
B0nVxy0JlfYhSVvNZo+6fvpe3KmzUkC4zE8lAHStyHGZR5/Q5Ht89LqGVpo+e8kUJHtJSpSMa0n6hSk+F9NUOCnvRwch6PruzqQUvUIBltWrRx+kkf3ZaJGdsTG5SF3B
ndkbChFNnAtJ8jqY2R65KuqEXCsBgq2TA0YDRx/RJHiKAhkLRxvDSz2g5a8WJYk2mNgAUH3vl5dYh901Ay2azFmmRXPNP9Sk+c33j4JcOELmit8u0i3JQpiiazWuebK/
Z5PdRw7Zzxq6USv9weJm2j/OnLSXQ09RcvTXUryAawGbPHvIjiIERCJI1GH5BP57DrB+nxNEvGHxGRqNMq88vz02+G5gXHeZTLUjRt+gs3yMtT5J1VYS6OgbfjHIYhEI
Jos+XVucqlYK3A7lrgmGNsoIWiKhhVe4oifNz/kLZLlYSpEmwgf0owJbN6E1/g/7WnZW9Zcs354QtM2UKzzboFDJC8G/JjUVUW6y/YgE+JCE3gtIYGDNgDcBqq8eNgMj
pK83xfIN/Qorawtbav7oy5MozW77ZaDjE7FpYZFAvkrHFy2p7qJaKLEluQ5Jj+IHyobrT+eirbHqrAUCDzElc/R6lFNN1bo50DX2fLfA1sMUg5N7fiXKoPiWu0+/EV9L
FrlmMs+go8VQvfRzYoQMLFD2Uf+NtRVoE1mSLpeekDHnK+ufgIt+iw47BJS/k5wC0+UB9Jb05vs58uL5+/uPvIWrEM6V5YI4X/i7VuWOc9aXBSx4GqDA0VSGr46p7Xuu
txJItiBWLRzR10wHmEedsLqQRIqCkiXDqZHfzU4e40/qQyRncurkRGnYc/E/NvGsGTCBzqc8dXwaIOCKMji+Rb1sKKi4Hilxk6qgeTpVwjBHRe+XNl10bTP6wQkvMNOz
CbDhS59YtTD5aLjVh4OzLM1C60jJ/8+cB58DYHmFYjnpXCH6Vj//RLUzHJMhxOwlyn0R9lG0muOQkL0IjABbNaaflA+wEaEjttrUOPK9SLRujGWmdtl6v9u4NJmfi6Rs
j5umR8iPbQaDi0evz1tendqCcCfng21wssCuxmGCFblMU5Lkq5Qc2dnBI92vVeeazOQl7I2D6nL/GU/Z7/TN8AtF0/nO/Ouapuugpma8YWhd6u2YCrhgQ9ywQAVv/cY6
YDGGpJII6+vHtH2hKaKVVI7L0BzDHH9q3bwAB+1HvFXiSqPxOkL7o1LZrkOLLOwbsP8upBUkuTpIYkASMzpTVSoMCFB+ono46v6efV+6Zf3r0cVGTNB9AiDhkxw2qLFQ
Q2Kqe9BVnd5lNURWNNe4Yhw13p6Z1b1TiuYgP61dDpP698AuEXkTxgzhDPGm3oktgzBSZOnMaGeLbnEIZ4w1Yk3ntRjeYtFU4+DcTLht6f/STGeObs7fK9H/zE6InBQ5
EcBwlLRKWIMn1y0N0RxomOpDJGdy6uREadhz8T828azdGI7rAmY9V4x7ribpmia6w68hJ5xZgz3vBr+7xtZmxw8br/PLI6iurdfG8iqLDcb7HhSOl0cfxLhlA7PYT+y/
nc2nythSHaDe6NZsUI8y2HPhh6ROCit3DtevBUWwMKBW47D3lJA7/VDt8o9h9AucePbKIiXIPqpWrgP/8SN+yW6MZaZ22Xq/27g0mZ+LpGztgAP7P5B2yLzF80YyXuNY
2oJwJ+eDbXCywK7GYYIVubT1PW7PcUdEST2STIdkcWImZq9onA0y+E5mLZHWxWaIYV7bIRLMQA1XbMwAa9Vp8iNVB5ECzBE9z1pTpgL7e9DgKLaEevjA9/ZANKSfQbd4
24J5kNShQ8Na7+idJH+EkJB/keYmgETpbFXygYEtO2rS5YM2duzTg2ukSGtmjyLTWhEeoCF3s0/bYRQKB/YkBumswLoqm6Sd6wokSY+txFx1N7oixlww7/W4L1Jg6scb
MLgHKWYFYRh4Y8KBJYA0rTN0F4YfXjIWOiTCPJ1RuP+5jnP9SIdSrCwe+Y6uV6lE+GGHNRE5nixUxLHuuDeALtJMZ45uzt8r0f/MToicFDm28HKkxb+GxvSuPbfmmFTa
CM2PFlJsMuRYhivYT8LyOKT6i/u4tLtozhXGhN9g28luMZ+8+tL1Jq3Z9j85eugaeyrESgKysKQ+pnzbnpxh8Ngf9dScuKe/kbbe3/GWUAqQ3U9q3FAufoBEPwYYR/v1
BFI1Q0d0N5VvTyMAewe9acJ4aVU78MKCa/37RhMQ4hPk2O3SFMSrbP/KQmg82T39L+QQZSoS/BYqTFTMzbEqF+KfC+7elZVTzlkW/FhjGlHagnAn54NtcLLArsZhghW5
l5b+EQFzOPy3GJbNo6v9ELceZaF2CY2rClUzoZfz/uWE3gtIYGDNgDcBqq8eNgMjIPqEVY7SabrpQ2qGRcwADkdsTxHSMe8UaREA9s/I8YHRvU89+rpnZ+OdUHpA/6ho
i5IpdFCcD+FVTbzsNb9+2W5fz6PfFL2v+jI0Mcubjy5Qh/AMBa7Wd0gIbPFL+XH5qXzMXAD1ZkTrDW552zGG1RI2XGrmVDhI/aHvfbK/P+yhHFWkq9+kuLEhimzpGnmx
dW8NaiGLZYI+nOr2eQo/pwssUtpMXFjvdawCkkQSK4U1u5kvp76CeOXEzyb6B3NI3tg36JZIjTN8D7VQ9R/VsjFXOjnuwpbGeefU2sloI4MIzY8WUmwy5FiGK9hPwvI4
XX7smQ1jJ8HZa42ZxQ/Ql37KGipBDnGnIX8o5QmthK8kWbNyqBzuMERfWLOuejlk+UyYw5BvbG+n7StJDW8Z0YvKvqUAxMn1Yx/4GLU9PJUWGLrFdMZUiyxfD9xJlDdf
VuOw95SQO/1Q7fKPYfQLnGSn0yy0ykwp18GsSaX2gAvMB+9cadiOnkTQ0lTocvF66rR1BgqgSWIjbsmijZxWSvXIkaNgSvgGkT3NvAYFid+fhJiYOMSCtk0VnFrGNBgx
/yHMipOGpg5J0c02dlICZypB02C2d3hVYEehXKvG/KwxPgfD6CP3ldraBVqF2ggkR2xPEdIx7xRpEQD2z8jxgfVeEx2OOfTkTEqZFv6Coz7KiCbRJr2HgYyrX3ljAm2I
ix5+UUvP/69jUT2Frv7VmRSDk3t+Jcqg+Ja7T78RX0tTdr5mhahzATLPZvBaU5Z+nORPN1l0bJpCG5eN6bImkSR7SUqUjGtJ+oUpPhfTVDjdYTa4Bcl0RmAP5IgFDZHl
rZY+XdSkH4lY6omSSWNTV2FerQeGniL/O5i65OkB2Mi7HMoXjBgX9ve/tbOcOUgj8vIS5gNADYeiybUG3GnU6fSp/0iSPsHvF4nQ6/uj8Y2AKv1oczoEhF7JC82/lOrH
A6EvQWzZXRgKAFppQ7PQTqRB9lyUJWWYvE6t2YNfuqRx6GKFF5jZP3QsndcvBquuHmI52bgb8MroS4E3rN49+ubIkRfuKFXQ6g0sDQfsFuNW47D3lJA7/VDt8o9h9Auc
Dq0LPJphanVmDUZwATVLg26MZaZ22Xq/27g0mZ+LpGzPKRFrFzQ3yGBavoCegn1J2oJwJ+eDbXCywK7GYYIVuQpEWnprnG9payQeShO+QE3HA8ngbntTFOvdKRUGrqF1
KkHTYLZ3eFVgR6Fcq8b8rPnd9Stpc19zddyuA80t1jtHbE8R0jHvFGkRAPbPyPGBvqWf7Ep2or9QKj0uOYhebYuSKXRQnA/hVU287DW/ftnB5tb7zY4+H2q4kEVQKF2F
KgwIUH6iejjq/p59X7pl/UlaVtui0uaLJPu4D53kFdIfNY8YDcaZ6T0tH9CrC5VbJqmt2xDuMq+x5eVLCIhvUBEA3v0/mPpVQV1xxwDNqBb1p78L3zb9NpqeLEVMWduF
lUzpRa2whPd+9Nh0IZbIsVEN0XFVS7qPH/APwydBTrF0BFtBoTSghIskonKnh19j6kMkZ3Lq5ERp2HPxPzbxrNRvlenEoO/Ce2v+Kb5/uKQDoS9BbNldGAoAWmlDs9BO
HTYNA9l4MxMSAyET+petKM9Ji9MPufYM/J7P3XKEBvPet2AzAdyznEcrFccO93DQ7WsthKs/K734r2p3LZZJA8J4aVU78MKCa/37RhMQ4hOQbsUn5n4E7jZSqb4elqF6
wa8GWQG04sLNezZio/fLvjS8lrkb1PUYfN1RvlxrQrIcVju+lWC2/+2wF6i36qzBp3UY30pu2dbYl4N6yfdEKqNkkrDT3sr9mnaMHDmTl8GE3gtIYGDNgDcBqq8eNgMj
sqoX2Ldvq3M3P/TwnKZ9RJMozW77ZaDjE7FpYZFAvkqpnIMT/fXVTrbWhAa4U0voyobrT+eirbHqrAUCDzElc39la8bZsH2yCkhgrkKyxIuShFEPum5NWjpCgqaDqsAB
Q2VQN36nGesojVLaFshcZR0He3RKeELPAopqrpBkvm0cNd6emdW9U4rmID+tXQ6TOZ57wD8G/xWK6j3iFlZvAK2WPl3UpB+JWOqJkkljU1demsdVfTE8kjv4X81L/lSe
0kxnjm7O3yvR/8xOiJwUOVJo6O2XZM1tkJ1wyy5hKW4IzY8WUmwy5FiGK9hPwvI4vWO/qkoi7cbcQEy16J0X+gOhL0Fs2V0YCgBaaUOz0E5e8rs98oyI6of1MIGoZe0z
lpkNgiW8alApkCzV018os/ZJLQqGCZsQM4skFfV66xKjWOwe+XO+0Z0hCiZb+v+hVuOw95SQO/1Q7fKPYfQLnBUzUsDY3Kt6PSI+tgc9q1pujGWmdtl6v9u4NJmfi6Rs
+yv25EbmiX2wiEkq+wPjmtqCcCfng21wssCuxmGCFbmswnorwIxcr8Jgu15nrbwGh5cxSyNSGLv0VAYLSIj/roTeC0hgYM2ANwGqrx42AyN+kod7mz3S9/r35ujF65qr
DT2KOrsT9gjx9wo9umnRPz43i2HwsdyN9HMBV1yZVMCLkil0UJwP4VVNvOw1v37ZXl6TcgJJ9DLFq2MuQO6U7yoMCFB+ono46v6efV+6Zf1nyjDvMGE6bXvwvn3khVEw
PNO9J8QnbN83KYC1ZJP7HakEO8NH6voRfuuAbpYKNce+OMr33W2mTvPpIxu5AIU7uY5z/UiHUqwsHvmOrlepRFSyEFwznVEmVuRn985uaS9RlWYNDnV6+Fn/2y6QofVP
TDuqbjKs1S6ud8HWNvsU0OpDJGdy6uREadhz8T828ax/HpkmFAhkLQ8mhIgXNkfEeZ4JQKk86JlFzsPZKQiIU4uRDNo/VO2gcFfQNL2f+PpNpj6FhGtdCMjyHQg/1Ss6
kN1PatxQLn6ARD8GGEf79YZoa6ALKYBAFQ06mSLFJ1XCeGlVO/DCgmv9+0YTEOITEp26BxmqH9TI65w3CHvjgsGvBlkBtOLCzXs2YqP3y753SEjD51PD3gfQzTXqYUzG
UpEJcA+JoTc5gSn25PctGLzJ0jzt3MKACKUWarZQGZjj4icNwqs7QozzLQjwzX2KMWJn/U374nmauItfuJWgXlHfv8Qa8dlCMFbnARS+1shHbE8R0jHvFGkRAPbPyPGB
EMjkehCn8/7ynkDR4feEC4uSKXRQnA/hVU287DW/ftkzSCBZGfC35T1q8ga2paY9gOUHl5mtU2FFNecuEZLm5eOLANBvykQMjSDiK2wIB64cZvfZ/vSoXixI4tjiHHMq
oRxVpKvfpLixIYps6Rp5sdYIZL5gpPo0nLM+++K+7cYLLFLaTFxY73WsApJEEiuFeyPsoMknGjnIRKZlLNiW1N7YN+iWSI0zfA+1UPUf1bICH3TNxPhrlLFp7WCNcB/A
CM2PFlJsMuRYhivYT8LyOA2BK0/9pNeO6+/qmSbQyM9uMZ+8+tL1Jq3Z9j85euga2nza8F6vaRMmvE9fO2h2wdw4oXHeVZUE/22B+MOuTVqQ3U9q3FAufoBEPwYYR/v1
/MBGtPvSDBi4OE9FtTDWzU+KPsnBYzS2ovnuXxWVg8/EYJSqT4/bYDVW7U0/qmXpqNEuuY5Djxbc3Je5gZMHOzT+soq1BezyWMZUnMp5Ojr1yJGjYEr4BpE9zbwGBYnf
Ymytl9Pw5cIpVM8DSNgtTHnOTSCOEtSM6DrCGI+Z6jfOJDnblkvrIXN+wYqxD/b+tpcp1RHvtudPtsN+W80vEGtVnLCh2Gg08fjPtfH7mm7DrCCH3O0tlGz7FYbIW034
yogm0Sa9h4GMq195YwJtiGvpsN+i52T23rJv8tGedAsqDAhQfqJ6OOr+nn1fumX9+6A3WO/YF1PbrloQ7W444RsoD+OWI+Of4OwDuNtlTXQke0lKlIxrSfqFKT4X01Q4
e1A3r6cSQgXiUCWt/NeIfQssUtpMXFjvdawCkkQSK4Xc/xiTUyipfGs75rUIlbJwUQ3RcVVLuo8f8A/DJ0FOsY20xegAoIbZ76Ip/xdVE2HqQyRncurkRGnYc/E/NvGs
ugyby2V0wunIUMIdgjaSz46r2Rf+YI0TQzTiqQ6js1LnV9EDXy8EFFW0U2D2680BXDWP5/eX5BCiFy500Exd9pDdT2rcUC5+gEQ/BhhH+/Wh/ThSBk5lsrY/2yEYqer5
T4o+ycFjNLai+e5fFZWDz3H9x1TiMzh2BSEeXum3cvnBrwZZAbTiws17NmKj98u+cgn6bXYeGMWn4gvNABiw5x5nBMwLT+sElcLlAqzq83DWMDmSwiPr9svxMeD32DMn
6N/6+xcUM2+WfRRi2qPMH+zzOnG81fWaUX2+9m5kxvdwR02QvK1n3zdOC/zIYICuDT2KOrsT9gjx9wo9umnRPy26HI/377r3P3EM2cJptdTmjYZGTPpx5fHkDH12aeTG
Wd09kE0oUfmgtpuZKuzvIyoMCFB+ono46v6efV+6Zf2rqwmqiP9P67OqoExLXS6DMoN5srP4tVRb/YN0MTNo+CPhLhIkQhok5xoz/wYVGYV3h2mqL7YyQflNs3xqEjec
IOG4W1aFTUfJefrZofanFhtNECmKULywqnY/lybvJzve2DfolkiNM3wPtVD1H9WyBt2lm3yPPaeUXI+HX/IHTwjNjxZSbDLkWIYr2E/C8jgJdxEykbKONnLPMSbs6GuA
aGT8Nf0pxMo3xvwe86o01mtfQXerXxA/M5ycVy88thACvbljE2rOP3GJ0vKJEdSGi8q+pQDEyfVjH/gYtT08lVPQ3f412paMlP/0pkT3AndW47D3lJA7/VDt8o9h9Auc
kOFVxEmgXpYS+fR03gFhx26MZaZ22Xq/27g0mZ+LpGw7os1WJxrFuWqqAh5v3RbZ2oJwJ+eDbXCywK7GYYIVuSgiuvyYuj0tP6qyhPsDnNe34FoOtrH4Uqde30x7rr6Q
hN4LSGBgzYA3AaqvHjYDIzXyylP/CFwjyyYzXEMIToGTKM1u+2Wg4xOxaWGRQL5KiAD3iQwtDLr9q/KNSF7wjsqIJtEmvYeBjKtfeWMCbYgHq853kiEbwPQL8QvamWOb
koRRD7puTVo6QoKmg6rAAcGSLXvht5MQVNalHoaDKtiagjuQbmafueO4r5cUuT2s7ggaiAbz4f9+gIaN35PQrstBtgOdTRS+SbDNbs6anfmtlj5d1KQfiVjqiZJJY1NX
eNBFSdycFsoPtCuMbD4wCNJMZ45uzt8r0f/MToicFDkmybuF+4vVKy+AeOcgWG1b9Kn/SJI+we8XidDr+6PxjXvt5P8j3xyAGxkRgF0qNNGOq9kX/mCNE0M04qkOo7NS
mPM58G2533ogkqCNOKSInTR/hkWo1a20+1LSxiMk9amQ3U9q3FAufoBEPwYYR/v1IP5JlTaAaojGziWpJy/R9MJ4aVU78MKCa/37RhMQ4hM3sR++BFjnBxuUejDwv5ye
wa8GWQG04sLNezZio/fLvsd4uxw2glezcWoOzxhSS4r1yJGjYEr4BpE9zbwGBYnfzuxzlHQBPgQzUgHZkHDiGHSoG8GZ2OdpK5mcpI+zJZkxYmf9TfvieZq4i1+4laBe
2rECaZr5hI2Kk9FpdzXr6ULZJnxFLR+05+2wLmZ9l/tCxkSz3Jm8JTUvkuSAvbUSyobrT+eirbHqrAUCDzElc8363CWPsQ0KZeVoxVzVO+8Ug5N7fiXKoPiWu0+/EV9L
ugv+4oGLgF8T7CE6JydUD5Y0GUWXT4+/GtH5v5q64EadmN5q3UQxV8RgxBZvKT4rromebQDRoL9m2nekvbnzEgssUtpMXFjvdawCkkQSK4VfKlPPVh0kh1al+h9lhkvx
3tg36JZIjTN8D7VQ9R/VssBMEzUf5/pgKG+x2BtBm87j2KSvYoMebAYY6iiN7r3PtEG5NtYxC8J1ciYuSnA8P46r2Rf+YI0TQzTiqQ6js1JpxscUakI82ZKIEyrEzxnZ
ENIl5M/YGhr7JANKrV4prYvKvqUAxMn1Yx/4GLU9PJVlKKX+eJm7QB99xbV4tdL3VuOw95SQO/1Q7fKPYfQLnGdeNKkQkJ/kxRStU5xvQtzBrwZZAbTiws17NmKj98u+
edBWmngDwGqFkE7beuJapTxQogrHIgddBkz/1N+H8D3p1xt8VIUzpFIoGCbqC1SbLY3nv7rcr6yROcm810oT1zFiZ/1N++J5mriLX7iVoF4n5AlmG4cGikxx0I4erqaX
R2xPEdIx7xRpEQD2z8jxgbhOLGw8xMY5TCZrYMZ9PZ2Lkil0UJwP4VVNvOw1v37Z0/Xi4aEMMna3uIHMQ5q1iVoRHqAhd7NP22EUCgf2JAbuqH/8xEmWKnPcuBRjtRbq
oI7SPLSyD0SYN5pP4klUvqEcVaSr36S4sSGKbOkaebFV8n0GRdOWb53Rc/7we0bMCyxS2kxcWO91rAKSRBIrhU76KHq7Wlp3Rejs39iuBbfe2DfolkiNM3wPtVD1H9Wy
ajjfZztGZpjT3Jfte0eWH+PYpK9igx5sBhjqKI3uvc+cZsPBZPulOUmWNQqglacajqvZF/5gjRNDNOKpDqOzUhoJH/AI8k0zp5GQneLjmbjViwK8nqs8Cd7/RY5hfL5i
knVfFikngIHMkgsguEwex2RZKzPf3bm9q8HIhlwLb8xPij7JwWM0tqL57l8VlYPPtaUC3f/GkUBrO0j6o84JUsGvBlkBtOLCzXs2YqP3y765bj7nSGg1JbV3CCU+uKly
9ciRo2BK+AaRPc28BgWJ39yEkcJzuvns3HWuluKiaL7saEu9zlujTV9nm8uKiT2V7PM6cbzV9ZpRfb72bmTG98quLs+bT3GTlA1x4FW6XK0NPYo6uxP2CPH3Cj26adE/
OaVkUM8lp1d79z69G8ZLk4uSKXRQnA/hVU287DW/ftnYg+jyouY3lwWFX2ZvZKv3FIOTe34lyqD4lrtPvxFfS1yM89OaAa6cUMk8HoezCDucEG3pFiNTT9QRfS5Vo+OQ
JHtJSpSMa0n6hSk+F9NUOEw5bFYnq4f91jkXb+j2/loLLFLaTFxY73WsApJEEiuFvWLxDRcaTMIiR9HhFFQh8FEN0XFVS7qPH/APwydBTrFcJgxsuzvJ6qPOjQTYyVmD
6kMkZ3Lq5ERp2HPxPzbxrMm7DYcDvbHgX+mTVcpigk+9iNNXYivKmafiH57yf2mYmtsRq6c3hrcBR+pPwX1MBQXcV5aT7z71fTexoTKu3C6Q3U9q3FAufoBEPwYYR/v1
EsrXQIErIKhpeheb4p+aqQ+00DbFPYUhGYk/d6t/HOJOZYq6S4kWW1OciPBaNqHhhN4LSGBgzYA3AaqvHjYDI7fPxKT1Su3mtzmD/rBGaPqL+g/CjMCBDu9w4b8c8UrE
8TMJwksAznUewo5SS0shI8Mfv3eZWtGqIFS/QZU8bpcghk77gDsK+J8sjd86MEKEIPkgf2FkH4S9fJig1YoE02iW2aPjjE+jCTfqKuosHMVw2jHPu/hM3Hn3++S6RlYr
ldwqoSC8L3+59ga/8M43wEoNnL1knsWEosbw0HzjS6udG1L/b/036JIZnsFu+xX79XWsKibcS5nY/m4SrvqLspOj0sL/ZNYUy8KmqBgnFsGLyr6lAMTJ9WMf+Bi1PTyV
J0PHRKLr87gjv2y87FFHihu2xEUJZvrUzN/yVAaZjDTT+Joq8hsNUTRUW0W4bmsAviQhwO5+bPWFrBb84YenOVbjsPeUkDv9UO3yj2H0C5y3QWp5AcdmDTlfypdUSWjb
oqdP/GXC5YT7gAdr5bI/HSt4yzJRwMwbtPp+vPYF5BGLeb+yBH+aIcPdCFvo3SLsDhqPSVAgQKTqmGzzjmtrzrscyheMGBf297+1s5w5SCMf7XVglqVwN6S2bpfPF2oq
DhqPSVAgQKTqmGzzjmtrzt7YN+iWSI0zfA+1UPUf1bJMjutGtjgaTHGej6+mDboUHDweC+c6YsqaWVt+FNO7MXMXdf/x26kWx7gAA2fjwJxlGOHwi0AQCt4rzAZWTf1D
R2xPEdIx7xRpEQD2z8jxgUdC77TRMUe3i5a+w+m4cH3xmYc0yOGILcC9MNYZAQHXyogm0Sa9h4GMq195YwJtiCdZMXEZMcSwUbCZojnD5p5Rp3rrdmUV+STh5+c7fGJx
i8q+pQDEyfVjH/gYtT08lRP+bwao0odhD513MIOpN0SE3gtIYGDNgDcBqq8eNgMjDppQIEwKE16lQnA7wfuLdVPwOFf40lQ2LzLJqN8XWhT5SuGiN/sQWS+uv7OtELhm
tya4cXpSTWb9AAzVx6088ShUcgoxtL5qmxVnrMJ7+6bfTGQmVTAc1WWBgJa/S+Bh9Kn/SJI+we8XidDr+6PxjTlCf+SKQmwiO73cVfez6pLW9Bejxq1SNOvKy6BCSWv+
IOG4W1aFTUfJefrZofanFmdWjGi78idoW9uXhbVLjT9wVl9dJa8j6cYpWlx9x7yCNSLRsClhvi0Wlsz4PRSlvCDhuFtWhU1HyXn62aH2pxbKhgK3gdmx8tfAunuOyjUZ
L+QQZSoS/BYqTFTMzbEqF2O2sdOY9iErg5RMU3loXtZJI2fAV4xAX6olsnZnA4jskN1PatxQLn6ARD8GGEf79cmcVpN9qRoYxoPdNVCHK7F4iPC91OPYYBbkvarYuc9R
E2K/C4B7FU9YI2/LvINQTd63YDMB3LOcRysVxw73cNA8yaZpvkGdMatQjvtkDAizyogm0Sa9h4GMq195YwJtiG4FEjwB6cNHcOppc9dxW0NGDshDKawXcd1T9rYdS9aT
vW8bCb0YY/2VofyvieOuBZc/95qi0KwrsVFHlvncGletlj5d1KQfiVjqiZJJY1NXGrSrhgMOUBHs3/o6HvuguHyIhon/bARRSEkjIyBlXWgPoV0S1mwSSPO/WySR6XGa
1I7GJZtbWV4clpn6obQnP6ZsQlc6hMOyV8pi5UDQnlR01VwkYPekZ5/kq7IepaH8RQeZghvvbzto2QWmwvOUnZPT6XgjaXP8DW7N0L6cbim7HMoXjBgX9ve/tbOcOUgj
md+qH/KW7xV32X3zKg8+hloRHqAhd7NP22EUCgf2JAa2OVC6CjsDgqzq9bCcsi0y8xtLAzE+yQTttxNZS+FR/PH2JSp9apZXlE6EcdGvhbJEx7SDuyF0S5IAc1wGiFcJ
AlDsx3bnBKZWACMZk303rgMtM3gzSwK6ngXDa/iJiZfFPs11Di6DXZPqxVpk0THsWE6IXobfjdUsQ1kvCfQkjSDhuFtWhU1HyXn62aH2pxa/4dHXFeCxJ0GhiQ8PvdiX
lf3UyQiLv+DDijxgm7dOjrscyheMGBf297+1s5w5SCNOhzY5nDCL8vcmFpUUsNkcWhEeoCF3s0/bYRQKB/YkBm+ZNrBrs21J6STrJBWnxnpZIrZHcqR2WYTYCsjpuH4K
kN1PatxQLn6ARD8GGEf79V7H3HynToB7pvhhOF/n8f4gP9yemTXX4gP2iKo6GS82R2xPEdIx7xRpEQD2z8jxgcEnVrgMuPK3P74C8a9syg4V5Tij+hYJ4pIxW16cJAJ1
yogm0Sa9h4GMq195YwJtiMJDhv5a4qiG2Le7vLHvLYQqQdNgtnd4VWBHoVyrxvysbDrrzjc/ThwHdniJGDLDlciZGu0YKI5ZOnB798eTkhwtzYmOMBL8Dy+Rf8imCddO
wnRsorDKkwOgMpc69Gu4i0x/sAE3b/DMH2sTPF8xmQze2DfolkiNM3wPtVD1H9WyidxZhdA/LeN3vx9HQUYI7JKFhgKvr6/lN1gqYBx1Kp6Q3U9q3FAufoBEPwYYR/v1
ygcGANInyIQx4KV8lTkiclcih5iD4p62FLhDPqVXTVWJX+l0cKldr9TX1cELIA+y/yn1++pKwdyClaaFiLdpuI1quJz5Qp751+qfHkUihc4v5BBlKhL8FipMVMzNsSoX
EtIqpLI4v3xnlScBAWl77wW7OQ93GCpxKsYB+PPnstvoN+QiaXfHlsBrwIZT5n3NYJhE2MOdJrcQeJs8otOojpMozW77ZaDjE7FpYZFAvkrhFAmSoXJJqyusb/5A4pFI
3CNjfUrdgcM5K2UCjUOiulEN0XFVS7qPH/APwydBTrHDGYLGk5MNho++S38yYRyYXI7QO43GDLuoJYYY4FK+xPkXSOoGL9CxHq1uebk+8IBMI0bK7gOU1wOZlAQETQa/
5m8EgvDVCUPWt4NAuFhhJQJWrEqDNg/EBgrRwZhhUCqCbPAttmy9D9+PdiuYODf6kyjNbvtloOMTsWlhkUC+SkQ8p/ec6nWXz48JCEoWEljCeGlVO/DCgmv9+0YTEOIT
i/zMH3OqSGskSdwugxx72NAEKX3dapJa2dkSW8FRFPEHMqQAUS+ZvRZFk4PLMf260MXhfKGXcnNdvTFTGhGPjvEzCcJLAM51HsKOUktLISOInhUZsyZ+5/FQahXFEWU8
FCRwycSN25sVqqg0I/0/Ji3NiY4wEvwPL5F/yKYJ106ZQHp346OhDsCYQXQdmO3c5ABDjeu/VOScFTmcHI8nGaZsQlc6hMOyV8pi5UDQnlQOaISmFKtmOKW5iYfvMg6h
8ZTNuiAncRlkxBoUqOYt8ySNhjgqldhX+sl30RQ/aJooVHIKMbS+apsVZ6zCe/um+Rx9oNX7jDeGNSuQ5AfXFXpBdfRN5/hMUv563Dt7aWkb4TZnTyMXZ4xqUhel9u5H
3rdgMwHcs5xHKxXHDvdw0I5UzyOcYzJWglVOtsb3wTu7HMoXjBgX9ve/tbOcOUgj2Fkiml8ZKqqfdUVICb9KAfYsBGgq9P1kEP9CAnQKdmOLdXeeA9HEaKczwrGyLzzb
i8q+pQDEyfVjH/gYtT08lUzG61RkUIhqfTl+DvIMhWaJgkiQiDjleQvzmXgdB56/G50xSk68S+Jf6kO82xsWSUCaAmH+J+vQGO0CVve1Pu6TKM1u+2Wg4xOxaWGRQL5K
9f7Sh6DfdznYHbRpC7ARqkdsTxHSMe8UaREA9s/I8YHfCJXhJUyG/P690xe+fkOX6bqsVpwlJQ1w03IUMzcha6SdHrLs/GOO/xbDlMZtEzmIbo6Mhah8FCquoiMKRB+y
CwhTJK6j5d5Mj//HI6zEGFewDOCe8DENiRjN3jJX8LUxh1VXPfaGN2G3kz59gmASujzlUzOzKTHqttRcS3kIvit4yzJRwMwbtPp+vPYF5BFKoLRaD8H1znV+6vbwZJoO
RQeZghvvbzto2QWmwvOUndXxRPfPzmU4H10kujzZBSXCeGlVO/DCgmv9+0YTEOIT3f3VT96FBXG7tLrmXs8J5cZJH1FpY56ut1YF0AMGBJcrp7//YemKTzBqgaj/rpTg
wnhpVTvwwoJr/ftGExDiE7dBankBx2YNOV/Kl1RJaNuj7Pq5dREJbZ7gZ2xtk5QLR2xPEdIx7xRpEQD2z8jxgd7XLf659YxvhFEGLROKCFZykImh/4G9fsQ/rRXUEiwe
ZNMlP18cM3JnVQq0QqdDxLbYfOn9u/HnGp3rK1Z6Nxm9+iIhGfe3ct4hZ2mAhhNMwNdZ66Aj/VNStCaDIQNljrbYfOn9u/HnGp3rK1Z6NxmTRsz3/8torEEsrmNuez80
SigKxBwgKVutx3YyNlNE5/vjo4/+pDm3lNTRAixVJEJqiyAmVT+ogggVRRY7cjFRcqn93w9ER0KY/W0UeRByP8qG60/noq2x6qwFAg8xJXOEBkVMe9IaKpaxcFRPpXAp
yobrT+eirbHqrAUCDzElcw6Id5PA679KYILnduvAxILKiCbRJr2HgYyrX3ljAm2IBJYFnQUZtKidU0idOPKh/+LV1r3av3hVOEoKPDeUKAspjvxvDjbESAEH12N4m7C2
6BMblUF6bulCH1xJf2olN/EzCcJLAM51HsKOUktLISOMuXjg/q+8ahPA+LASBWR6Rg7IQymsF3HdU/a2HUvWk0mUgCxpWYPbbZs+0fwbUt2keISObnxVrAl7QVX5zOTR
wnhpVTvwwoJr/ftGExDiE54fR0HADaqkaDgj/s3fJC+Q3U9q3FAufoBEPwYYR/v1/oIwsXzpWON9aWOv56Fc5oTffNpkVphgnbClFC1aGmlsrhXQSpj1lrLY4BmBLvnx
Y94XIU0Y2HdZlqnzpCIV2TByYh4j2JoYSEWvzvcdUnT52PkMn0dQmZvvkTL7e+gGGULQoS9YYip1ZYoS1bHZouizlcsHbJOFaOQyzbcsDYHox4iojIETWrNRBvNXfTj3
jWVTPVvEn+FFqJP0DHjqWAUDhEeJCouZIysnIebzDA0n+yxspKLqzKPcnzzxlyLwW3NpNQ/gFg0nc8y7UHfn+H76s4zk/99nkpG8k1oS0PQlenRwpnYlgX1Zj0RNEMPJ
9Ohabb91qkMmoacoLXMcc22mXO2wS4s967vhP6jo0q4s+F7mu17uP/jRgWsyx7FQhN4LSGBgzYA3AaqvHjYDI6KoCaIO4AvOA6zHc1Y9x95A6G4SPNJ8WeJV7nwQo6EZ
6kMkZ3Lq5ERp2HPxPzbxrHTHut0MQ1pRs5qVEQprKJFy8Kl5DZOqiMQwh4sg3kLTFNEg1sSa+4ePVAMrZSyRyLscyheMGBf297+1s5w5SCPrMVx3K5hU1cxJ6UTxlH8k
ZNlr1o3MznUQFsferIovIvb8fMdni17mHOQ/yISmuvjet2AzAdyznEcrFccO93DQkVqnKMM06Z369DSawodTC97YN+iWSI0zfA+1UPUf1bJo1fRhV1yS4ULvK7eSirg/
tCNfowHW2Ihus8d/rcha7sqIJtEmvYeBjKtfeWMCbYhaRFdsNdmeFU4QgrN/oHmyk5YprFIzIfhEwA4t+4z90WwaxmqyRKB05h3pXjQ2ZQhOzA+sJHh/DjUlH0WVMzyl
6TIKK4bwZ8i8OBeCm+6seL1sKKi4Hilxk6qgeTpVwjDuCBqIBvPh/36Aho3fk9CuVJsoNFdn9w8kb1eCApY2CChUcgoxtL5qmxVnrMJ7+6ZjH2xGim6nMJ3VZFxp6G+l
9iwEaCr0/WQQ/0ICdAp2YxWsSDafXfYqR/1Fb3gieBGLyr6lAMTJ9WMf+Bi1PTyVv0cPT3m/toPpHKsaPoNlb7scyheMGBf297+1s5w5SCO3t9cDb/no8F9drNhrOWiA
eQI0zeHzTg+xkt9lrbgsVfjmQxvrNX447AOWfyI0uZVHbE8R0jHvFGkRAPbPyPGBl5MEyLo9SrPoKZjddV94mzf+dUpp7dKjH6BCNWXq8oXKiCbRJr2HgYyrX3ljAm2I
FKOxvnnqbG57OJGtpq57Atd96RZIBR5rRzIEAgl+i/XT+Joq8hsNUTRUW0W4bmsAvbsCB/GsFE/k6iAfV+n25cJ4aVU78MKCa/37RhMQ4hNwmm+3VuHwfpmJV2j/8iVf
9SL/HazdyuUFoq1AnTngWBBRKwS5XGZFfqbS00K/NNiAcwAwp6T4rn5yK3d60Efv9Kn/SJI+we8XidDr+6PxjYplJsvecHlh7mGmjrZc0GSX6Z2CLLu61AGpCpHFcyYd
06i6DAolBJZgJmA7tmLVFPkXSOoGL9CxHq1uebk+8IDWKvY1beZSLBT9msAvQ9/GZ6WEot0jED0pGAnbEbm8nK6OyH6/VYggpG25RiJisezqvNJC6Q2cYuds5BmljXJC
Ay0zeDNLArqeBcNr+ImJl3takBGYxIhUo2TU4JhVB0TD/mjCsfl1Ed1GF7/bdQeZrZY+XdSkH4lY6omSSWNTV0tNweFlkPyF4ih1t8sBF/jKiCbRJr2HgYyrX3ljAm2I
D/BVuDCKRf3u9ljTfWduuF7rlAZryZYRQyI7Xf4JezVOxirikV2NQ3bCKYUJRta0i0vRXByjYi01joJwJWb1hMqIJtEmvYeBjKtfeWMCbYjY15v3WXSGe8FHSmwwDq1m
jcGQEyb82qidiiZrYcxiEMqIJtEmvYeBjKtfeWMCbYi0gRFzuAEGAo0W3BzHzISkxwfFhKpYA6PzIsb9tNKo5fSp/0iSPsHvF4nQ6/uj8Y3B9C4HpdoQWWD53OHIYn8w
/iwDQ4W3nUc73+65UbJB+ezzOnG81fWaUX2+9m5kxvcaoB5K4vnOJo6qHvWO2xw4K3jLMlHAzBu0+n689gXkEQzheFdXN8u0sOty2AXpytj0qf9Ikj7B7xeJ0Ov7o/GN
ojXjs9C0zWDFs8IeFwhsb+qGu9HVwCQ6COusJ79bh53s8zpxvNX1mlF9vvZuZMb3rscMcWwLU6NvEMNSqoz6+CfZcsbr8AS0IXcujMUDRieBmPeB57Cn0px+nG4PWjr8
fwlyLc962xAIiwmskKl5s/Amra3Rzvayevz313Gw3AUVs4AXo9k2KWI/pwWjShmLyogm0Sa9h4GMq195YwJtiAIsR6OhfAn+9OcTEIAVUomB/mSnUv7ovXZ04IeYQwc9
NuvgfdKgCYNLuWAhAG2VoskQpPO6i+67PVnNBSaBd1dqFlnOHtlZS/HROug4r7LyA94Zyqf9REzG3RXdUDRDR831EXv7QNtInYUOxgOd/8p0bgcSRZC/5n/WntOUCz+3
JATU+VnTpQdxaDsQik+z9Tkko8HdCdrJOIhYZmBqnXHhiDQ1aj3aqMC3ZpERT8Kce/VOffiHCWsZZ5M5pZG81fYyw/lbF7mxI4fRwJcw9FXe2DfolkiNM3wPtVD1H9Wy
H+11YJalcDektm6XzxdqKgdDlGPHxXEWJ3Uo8YISL/Kae+Pk7D3Cyn5N5tqNVH2iBqnb6l8gcqA859pthk4LIx2txOv9uoEB8oRhG/ahhxWdx/Jg13bl656shDksb9Lu
Y/uIKlARMO2nakeHfDYae62WPl3UpB+JWOqJkkljU1eap2C9BwvUmEsOhSlJYdPrEZKDGMPpWNXd1O3xvWcTdcuID2/3HLxDxvHdQWa/DXbolfSZrKg7TMUJ0mTMM5Od
yogm0Sa9h4GMq195YwJtiBajXJtD48lErnUdIYSFoKNSQYwa5zeKbKeVTK70RyEcy4gPb/ccvEPG8d1BZr8NdgXW1qHN5v6ml8kOHjroPWStlj5d1KQfiVjqiZJJY1NX
kQ1GJVCZ7AZeiFWk4YgIeRTaqYO+gYOVq7GIcDbwICxFB5mCG+9vO2jZBabC85Sd1mBfX8k2cfEguHYQoxhVN1Gi8K+QXQ+b0ucrpT9/ntO6h+pOLDrnMrx9Os/xOxmj
yogm0Sa9h4GMq195YwJtiI2o54Ebdky22pj+0z1RHFvj2KSvYoMebAYY6iiN7r3Pi+JxUSUTpyGxMJAnvxbKQh5nBMwLT+sElcLlAqzq83AOcl6+U41OcrgR892xdOhv
/yn1++pKwdyClaaFiLdpuLo85VMzsykx6rbUXEt5CL4reMsyUcDMG7T6frz2BeQR7f326N+m0RGQ6B4xZjwbiD7oQTe0uF9GysgupuK51Msdg5sWs3VWEa5vGnpFF61c
xkkfUWljnq63VgXQAwYEl+ihk73jj9UKXb1gGnRkndQn2XLG6/AEtCF3LozFA0YnzAvgoirw4yxlRcOMOcNYCz7oQTe0uF9GysgupuK51Mtmm49errq/zBFiD3R3SpQ0
e2zvzhUa/0qKhPZdiBUfQYUCORVWObNYYaPf9wBNj2NP8dMd/3OIsqOUcAocWq7bHUHpn9b5TIHubZSMliPraZ1gIlY0/EpYETXxR6OleMy9bxsJvRhj/ZWh/K+J464F
Mvkd3XE+76NAukNXzey9mYDWT46gIvUPwnr3wF+fa8A9FMJguPrOTK8Rc2O/d53PkpFEAHvAxIcZJQskbG/0ViEzBlUlrkU+LF+IfhGL4dnKiCbRJr2HgYyrX3ljAm2I
1MArccl4XYOVs+pj/0VmwqqB2gb3Kqy+/u7EzdDGgs3CeGlVO/DCgmv9+0YTEOITlVWqfvfDXxzTfsD/6zDhY3dty/Ot6mmZKBqJvUPKxe+3i2idn+4+yAXWCD9twfyr
lVWqfvfDXxzTfsD/6zDhY6nVjfLhnKw6f8VDjzk/VBVRovCvkF0Pm9LnK6U/f57T6g+Zy4yXt6clIeJYYj8cy1TZPGEdgHs+HcP/07zqnEytlj5d1KQfiVjqiZJJY1NX
6g+Zy4yXt6clIeJYYj8cyyq5jG/Rmy0NQDW3hDb0Eoitlj5d1KQfiVjqiZJJY1NX6g+Zy4yXt6clIeJYYj8cyxrobDxFKYLJfaxQzDqpmwJ/gxLMiS+gsr+eq5ub5cwy
ZcFZF4eX9X4du650aJrWvNpF5g6+kBABAL2rZHl+5rqm5OiLQ1cFMNPqd172kK6CRQeZghvvbzto2QWmwvOUnTMdqnTHEoS5ecYZtvj72r2mmxu+3BJENG1XVjzuwOTv
3A/PxgQYWgYJCytdn1VqUY1dmbJTdn5xFqDltKKOBK4t6Gj3PU3Pg9Cgv27+2+Uxyogm0Sa9h4GMq195YwJtiGguChAH+2iJUeWEM/XnhVzB5vSE6maHbz+09pht/oe4
UaLwr5BdD5vS5yulP3+e04M50MLz0x6at2bBS0CpAdnVlTFeQy/Wv1bpqYplmg05/eALy2dF3DC12Br9RObWR4hujoyFqHwUKq6iIwpEH7Lz5HSrtbg6gOfBSLxlfgqq
W4w66FnzKSZ6ZcGHXe1F5SmO/G8ONsRIAQfXY3ibsLb7fYQ0XuIYHzWN5G8fqdEhFgdpXg2y3LzfPvcfHmZe7y3NiY4wEvwPL5F/yKYJ1057b5lF3FiXolRj20JN3yXY
LyDyASmEMk/41Bfmd9wsI/EzCcJLAM51HsKOUktLISPsHeA2LCZg8gzb7/Cs8+MDxJvPb1YR97bsv3l54WbpbsqIJtEmvYeBjKtfeWMCbYhoLgoQB/toiVHlhDP154Vc
ExXgN8IkXOMibQzvq0t5Jd7YN+iWSI0zfA+1UPUf1bLnlBo9ErEpfMIL7KUEMeXkhU6E94g7mNy+accyoDIu9ZTEBloKbv+n5kG97lGqHDymbEJXOoTDslfKYuVA0J5U
y1jPIUmezd9DZe8Y5m6aSO5ioLssXWsOk+sHFXKX80hsGsZqskSgdOYd6V40NmUIVvA6oIUoj8GkSnRkfHF1xaabG77cEkQ0bVdWPO7A5O/xMwnCSwDOdR7CjlJLSyEj
7B3gNiwmYPIM2+/wrPPjA+UMZXjoE/P9k0oNvr0iDCLKiCbRJr2HgYyrX3ljAm2IeT2/yUl6OFdMQ8D3TJxLIcHm9ITqZodvP7T2mG3+h7itlj5d1KQfiVjqiZJJY1NX
p+5jzd59728a4fUek8rlEAj4ohy+IVYsNXTkK/8khEbuU1xXqfNcfYZTC0r3YbEbG+g//CI7tSCYj62FAXs62bs6q3D8K+Hd4QqUQte4PlExveZDShjZ1uuOEcaRp3AI
tth86f278ecanesrVno3GQEAbcHdD3ZcDXxrp5qYoeULQeYr6/UJxZeUX0KAU4VHtth86f278ecanesrVno3GQEAbcHdD3ZcDXxrp5qYoeW0qK7x8ns8AiF/wDEH+TTk
pRnrBbYW8cwbNg7Be/4ZF7746UuIWXZ++74xqR6oYmuNM//v+JdscnvNRQX8dKlVpRnrBbYW8cwbNg7Be/4ZF7746UuIWXZ++74xqR6oYmuyu0p2Stocct6bEWc5f9O0
pRnrBbYW8cwbNg7Be/4ZF7746UuIWXZ++74xqR6oYmvMGKPpn0ENERps4NwNI9ScR2xPEdIx7xRpEQD2z8jxgYrLThC32HXT7kEVX69UyAGVjjuaZWD2fSc7HI/RT02G
kN1PatxQLn6ARD8GGEf79cLpPBu33Sacsv3NyXdI1c7vKR+2yuc2PpaocpvCd7i3KkHTYLZ3eFVgR6Fcq8b8rKaV0Mkc1yz/zj3T91hXhdT478nJ331D6vtUrxVTgQEQ
SIca6qBaXyU1PliALg0zPLegm7moTKO2YiGDGSdqHEwy+R3dcT7vo0C6Q1fN7L2ZOmjYWVV0p4/2DgaDEpQc5vvjo4/+pDm3lNTRAixVJEJhKRmh/hBb114zswOPouJ2
UDJT+p35cTgDfuH27ebos1Gi8K+QXQ+b0ucrpT9/ntOuCyUSYrpDStbtXEOJymrRvmb1ladDvcyEq4a5t03B0A2e0iGxjyFcO8uQIvY6qRSSQca/OoZZ/ueOLeFn/QXw
PXcw0gFL+x0I8QAN2OIrD63mEPCKhtJBIzL3vNhjfSgD3hnKp/1ETMbdFd1QNENHcLV3vWubh6rtdWi6+DBlroJ1PacwgoLvn+oq/LGQwUzKiCbRJr2HgYyrX3ljAm2I
7r/MHQzFg7ErUSfLgHrs5tRJx/rtdbKB4Gcl4+omcYBHbE8R0jHvFGkRAPbPyPGBKMd1TcvnaWFRDGWMwaWjxjNM/Pfwe17gc3bHlSZrxMoqQdNgtnd4VWBHoVyrxvys
HiXvcI4guY5gvR0W2cYnDAVjovR8B7ut9XF9+kQBKvgDcqfXV4Juxwv77TiV47Gq3tg36JZIjTN8D7VQ9R/VsqK2thRXLThPFCt8I6GwjenaiUvQjsukb2BRKMt9Lb8q
KkHTYLZ3eFVgR6Fcq8b8rB4l73COILmOYL0dFtnGJwxRFcjBKamuoO7zlVe8/PNsVNXhqwX6M7DCZyS+O1SwZF8H1ZgKYKVZbSbtinljn3JYecLFrhv6t98eHjnKs12B
OPaDY24Q8djjsLtUaAWfsLw7V87q48E3KSw/g7XpIXJszpcCZYT4Mf/Hsc83qOyXwaT+WmxXHuHCWffIYuNIkIJnEIud/FJo+z8qe6iVNbTKhutP56KtseqsBQIPMSVz
j1WDcLIXE9/qyBkZjKo5GhNyazgIvQyxHkd0qmu7JxzHbFr27zL/If1ymFzDLrvEfre+OnRAjFH9h12KooHjSKaZmfAgT8gysWXC4ysNfDJzCDOgPn5uCfww9AoxCFpm
vc9aBNYIf5ztH7rA2pMX2nxsu4kDD2FYVu2/Xll7t7VM1+UlBv7qTi75uV/u6YGDsNHsoLwJraF/3pfYulQTOTlrf2hXCVN1zEJbu2INdUzTma0401444/gjwFPXDxbs
kQdsUk/5jKNdL8uTVmDi2jesK2tUEjNs+B930VJvL/kvTT5WgXTSnWbhA+3hxo/G+lFIP+EjMSCfueYeMwbM3W+/LolJLKo4/wVJzjHm4rvCeGlVO/DCgmv9+0YTEOIT
Zuwx39vDciPIv2+YssY9HslpWlDZoogMs9JT8twbSKJwTKEb8aw9n+SH9tauQFUf+g95P7urU9dWfniP+g400iVXUdWe2MfIpxXgbIl8o/I6QuaBuc0CN8h14scto6uF
IpAieFkRou3K/IdoZvxZWMR5ysrwxQo31YYnDlgyz59ywqFp1c025kgziqbF5UVkbCAsLjLsTNY6Gvdq5TZRpevbMMISoai44sbYZ+T2+7XKiCbRJr2HgYyrX3ljAm2I
JryprLDsfWvjd9IOaMsRqKj3EvyHH4wgLZOyFJRlRfrJQQxoSwA/YRgLVshzbH0ukN1PatxQLn6ARD8GGEf79WDnY8gzlAvqocPkr5zHtB9fCXUahSeRrnsuRYNJ4h8A
Yu/qOZLbNgdQYvmfDw87vQEzNt/qntn2Ai9Lp7y/M4scu09gZlZiPM0NVkhATLxlucRFCxpdyQJNfj4S2VwAlNvt4t8BRHg+3Ex8qGvNZCd4IU+NIMx6ywyK2jWU8Wys
WTB3rx+PxwjPYe0jHqVblgsiFw38YG/M62rrg1PSyQqpWfmSFfMCG90dTAX1Ys5RK0IEM/x4Z/AmmiRaImznhSvI6jNkl4LMjTGt7WPrraMhcpYCGFn8n50xePkMR/o5
FtfQnl2O+fcS5sNiVocTL61kkEixcLBAlaF8qZu0P+s9fIwNoRhZn2rP25pfju/sCImtcA334jN6ckHyXoWGbZ4KqCc6nxAfdCeYEaTkzE4sEtv8KUDz8TWEb6EKeScN
GT2feqMfpyCdS6c3bjY4zwiJrXAN9+IzenJB8l6Fhm2eCqgnOp8QH3QnmBGk5MxOof+PR1hZ08HcKXeFWyt5YAssUtpMXFjvdawCkkQSK4UOkV/HcN2gD43JD+O1a6jq
hubch2BapsRhVJFV6YMH6n4vL0x+qaq6jNrpf+G+gQnH2HwKwmS7r37jODneANSNZcrFXxMfhnpVDLIKMAjeXCr/pysRRcgK+nqG1OAZUmc46yEpiM7rAvRjD9JE4Ncy
XhGf7mikKVef0telrq/m2i4CnyAETTwf7RIouEdoZpLntQ1Jse/lwgJ4ZxY9lwUx0ul1qyu+rszoxclaTKf0degFBd+ge5O2bw+GdPYIvB8FAtntXDDwHHgwesibATUs
57UNSbHv5cICeGcWPZcFMZy6Mwfufn6jd7thSQw7trfEoABEUiRCa76ggtifRCfjrGJoAtf65lHdxrKG/um9m1+2i8PY4VHDSetcGXJjGlkhlnmxlJX3519/lcMazP92
PhFY3JYZORjFTahqBzO6gqlZ+ZIV8wIb3R1MBfVizlENtiy7sL1IXvRQaqWEbssFlsHJublyYjZc2/OX0oUlROgFBd+ge5O2bw+GdPYIvB8FAtntXDDwHHgwesibATUs
2oygxcPbw4DaIr4fEU5qbTOJwdYJFKUkjH73w5lXLMTCeGlVO/DCgmv9+0YTEOITZuwx39vDciPIv2+YssY9HiPVevFhnOtv8vMzl5ZVWogHixpD36CLPtvYDiwOOOJi
ZcrFXxMfhnpVDLIKMAjeXCr/pysRRcgK+nqG1OAZUme8/dlxakEHoz9mV6f7W6nRDihf24kmvf30hmBVt9GuiyFylgIYWfyfnTF4+QxH+jmbHyT9yFWz97OSOS2+RGqy
RE+fkGkbqs7jS6K+MZMSB/xUHvS748xbBic8fD18R50FAtntXDDwHHgwesibATUs2oygxcPbw4DaIr4fEU5qbRz9CDWZThBIP40KPNI4WIvCeGlVO/DCgmv9+0YTEOIT
Zuwx39vDciPIv2+YssY9HlGmpLL6RBw8vONMWVpjMW1HbE8R0jHvFGkRAPbPyPGBZx17dNfebIKSP0z3pQYgSBhK/aOd1Z09aA/YTOn1Ol+Q3U9q3FAufoBEPwYYR/v1
ub71ftjGITaqYD7qXfX/jdE77xGdTUZBJp1FRGeeCwEjfF+n9g60zfMMDNBYuxweCNrmSqQsmtYkF/HIyj/c+Cr/pysRRcgK+nqG1OAZUmcZkowqj9WyMB2Ut1hedzMM
smq0zXCJisg0itRzPCYUpwLaAfycvrFA2wSsvHfrmxEq/6crEUXICvp6htTgGVJnphOSDvg52dDMjZqwHtb4l/hGb1ANrvK4+GgbM6stj5RRDdFxVUu6jx/wD8MnQU6x
qYdkhv01Bs3AfJi82yeYjHK2qqlj0pAerlEhy4+NG/1wpBEjOqfwSugDobh+Ikk4wnhpVTvwwoJr/ftGExDiE+p9ngir03FT1y6IRZ6wITJZbu2qyX5EZhX78DtUMzJO
FolCJRw9+WVfvRh03kclSQLaAfycvrFA2wSsvHfrmxEq/6crEUXICvp6htTgGVJnAsCcpEBj9i9LGT/ezIM7VH4fGntecJ8gaPJZHCB2Q+o4O8K5IX5RLEgO8pLa41bO
9ndtgQs0mZAJARlpR+WkxMJwq9YJdNHnGefyjnA3i/aQ3U9q3FAufoBEPwYYR/v1ub71ftjGITaqYD7qXfX/jZRBqRajFPAdeMDVRUom808rG3zeVhs9kPC5JozYtGtH
R2xPEdIx7xRpEQD2z8jxgShCIUlj681zCOZoMKzKIjiokTQU5lhwq+BHdlSN8yIJIne66wPSL5HqGpqfHnK/8wLaAfycvrFA2wSsvHfrmxEq/6crEUXICvp6htTgGVJn
6IaSiZFiqqUBYTuZd4evCwDpco8sf0PlSuLNIJr7x784O8K5IX5RLEgO8pLa41bO9ndtgQs0mZAJARlpR+WkxKIPPdgXKbiS1XCR40V19bzMR0sOE+LTX4h4bbavdCKW
X7aLw9jhUcNJ61wZcmMaWVJL2KNIoiftCBb3uCW0pO5w4hqa9MrI1iNiLDiL+RYRs9NCw+BmPDfPC3eBxNxpNJdE/SHeTk3F9kSdwal0JkGTKM1u+2Wg4xOxaWGRQL5K
KEIhSWPrzXMI5mgwrMoiOKZe1wkJ4+j4I3Jf68BLGicLnAGtOy6weyjgAd0MjOckcOIamvTKyNYjYiw4i/kWERY3p9vz9erKdGbuT9QeSB6d2pl/L5wNRkFN0khXyCOe
73ak/6ShZDl3FZJRwgDzZKnr/4n99EXyNTzBYPEI6HWT0mwGaq3YllErjRmt84H/uf4LZhlyXJftSMjby43Y0ovKvqUAxMn1Yx/4GLU9PJWTSnXYEL7/tQfdRt2rcwcI
k9JsBmqt2JZRK40ZrfOB/x0hTSu2L76HJm9+1IR+uMsyH3UQLN27/0MbVbwpAAVTbmQFGg9zTqlYjt+UEY1QOq2WPl3UpB+JWOqJkkljU1c/F+h2YGiZsQ1wYDnnuJJ+
q1mJ4gebghlMVLVwTwRmrkLZJnxFLR+05+2wLmZ9l/tjqpgmPHhYKix4lowM1RVIq8jlCdQn7IpIOp2efOrMQLGNH720jcdPjCanzY5qcElvdevExFH85W+mDseR5W5J
ShRO4KmzTpraim3jn5Id1ngKE5I1QJ+LyyJaLyzc6rXCeGlVO/DCgmv9+0YTEOITS0XXzcxsJWSF+hHl9qZcBUCEt1DAJbLt698th/KwtkK9j4b+2WyrQpbTopmuMgK6
lrvUkBHhgpZB83OSuXA8zzbsABwGJ0T+DzzIo75j3ZC0GRlqdPQdmujLIPvXfcoCyogm0Sa9h4GMq195YwJtiMjUHhGXhd56Uj7dAcFHjGW6joTJcg1+PGLloBmFw6B3
aPx7CCqD12UlA/I89e/F1mlSYAhpUerxTo3AbkffIv8I9t8Z3UyWilibXzTXvWNlShRO4KmzTpraim3jn5Id1te8xqsxP5bUwq3ipKZGauotEMnPrIBuwt+bx8yeZKYU
G585PVlNi2E9TosT0fmx3Dv/RYEUAICvmzC1lsP35uqYx2SPEuOcggAvrW7aTyDnkN1PatxQLn6ARD8GGEf79Yif+4BkvgbXG/ahWdxdrHLBVyJUfLZ9A5eQrXm7Khja
dYAE9ZcdD8R4w2TSv3aelLeLaJ2f7j7IBdYIP23B/KtGDySmfj8konTujqUk5wybO7GbmOgvypH06RYeriMWJ8qIJtEmvYeBjKtfeWMCbYjeM+J0ejbGcqPdj/cnxqhO
mUiYX2u5zHZ68S1HHf3l86MDh+XI5Yt+4QNTnWH+XL3gQAHRRhAoh3D01y+TnTA5FJlrJtrB3i+ShZmwhYuJex01tnl9e0vOFtNwar4LoSY712WCVXDEUzcr3vJN/M3r
LVfVHGiQKTJ+di0hKPRNr8XEmNO6XCg+2M1zKUoCa4xVm9QFYz0hJLvSVPqBA5zEuHBRsNPlgswwvQZ0isieVirT7RVGBzxUV1ob9UDhKJA9Umw8F/8vwg8lE/guR8TI
1gnlQ9vkKsNBFsP5W3pFPGe+hfUqc29f2xzsQvE4+kne2DfolkiNM3wPtVD1H9WyzCXduu7bb+Ug4VnEtEtOnnJI3dtYdEprvuilBeifbTmtlj5d1KQfiVjqiZJJY1NX
ilgyqZ3mRFNGnHD8FnlioKmuqQ2Ea9SBZNuMDRsBKu2SOgZJy6WDF2flx6tqCPcn+Qnewv8i7g3WdY15t/lAr+IePStPGhnptG5vwBOv6+YlmX5QGapzVhu6TIKm///8
Lci14gk57mLmrToS4XZbu+IePStPGhnptG5vwBOv6+YhaRmokyJHlfbNYJKtK3z+4Brcifyk7XoSu7SlKLlBtQ9599uYJgDHN/4piCTz92qmvS1HN3NmjK52oHu08mB0
38AgRzDvaFrNT3sFO1PikANgH/jDChfVYybm3yiVierKhutP56KtseqsBQIPMSVzCYz5N0mcSa1CzgmYXzPKsjX0UBDNPBneBNvKiSHfLFzOHFE6JzstY3YXRHigquGY
a74Ly22mjuoWgK8IrtyyaHbhXeSGUeqVHvp7GPz27DAy/Y2dBwqjfW7CknAL0Jsbfw7L3OlJXtAeZBNwTotiUosn/9Qcc0iD03ICXSv0JjM21edd5XN/3hBGKeSz/jQR
YOdjyDOUC+qhw+SvnMe0H6H3die4bKA138f7WaYmlaRu7d6pLk7sx5GvInnpt5uiqWIefSJnFi5o/LWTG0jsfNaKa+6wcNvIxDjX51kkaJr8PeeqZkOvyjq3Nat4e1CH
NBlX0T0Fb12NVKzc3NXgim83ctCJxYoSrRh4A6g99bx/72CUDJtBbs2/nMughw8dAlqp+8xjJ2FUOY6BDirKA5DdT2rcUC5+gEQ/BhhH+/Vg52PIM5QL6qHD5K+cx7Qf
2Cls5QF8YIw/djNn/W4e4cOEdeguBsLrJDQzP5+CO5ccu09gZlZiPM0NVkhATLxlC7gyyL2M43HR8ff9ltDfBmE5K5lrH7zIiFY+cEddSOVRDdFxVUu6jx/wD8MnQU6x
82w4EaX7DfQ9sOfGneP7itfrXR9SNqaFDoSCujoqd/iRw2ADD7DKV+ApTrRDJrYOa5HzhKj76hWYUSGBtGBmKgTXVAjlkaqkVydCznPCopjHpZeiF7KJkij9/uqIYwhm
R2xPEdIx7xRpEQD2z8jxgUiBxKlEj1Q+cLWn+44TkgfMB+9cadiOnkTQ0lTocvF6s/M8embq0NuYYo4hnuhp5Xgqx3aM+hqrL0pzF7H5GAZlW01aUONYhMCgq2Y6pcJ8
BQLZ7Vww8Bx4MHrImwE1LOLX2H2mXotc4Lr8rPuTVQctO4pddHQShAKyVbpnFZ++wnhpVTvwwoJr/ftGExDiE2bsMd/bw3IjyL9vmLLGPR4qwS2FouNsA5pH7iGc6a5X
mBMyk1zeVfAh/ev0PaMez2O6vTeNsR2iRaEOO3TlB8n5uIa89ITr6JGPeVedxgYM9RgASI7nFDgxbcwww+WyCNRJ8ePi0tWmzAItR7OXNGWsYmgC1/rmUd3Gsob+6b2b
/zowf9w+JeqKUpBd08q8IQtQpGDZ/wzR7a+i7EOPeXyw0eygvAmtoX/el9i6VBM5OWt/aFcJU3XMQlu7Yg11TNOZrTjTXjjj+CPAU9cPFuzGG4a3YqCnznXqa1DtowVV
rV4lKp/iSh96LNHj0oCfi6liHn0iZxYuaPy1kxtI7HzWimvusHDbyMQ41+dZJGiarbfBfAyCZDBZdVbipSwI88k3Ac9DEOM1PMVoswHMCDepWfmSFfMCG90dTAX1Ys5R
dbIlxKcnuwUd/a0q3jTA1RhsgfLdGZ8DvT66CNcMeTriHj0rTxoZ6bRub8ATr+vmZx17dNfebIKSP0z3pQYgSNwlF27qDMw+hIGgfrBWkslJhQPtzxprb7n3SQESUEI/
yogm0Sa9h4GMq195YwJtiCa8qayw7H1r43fSDmjLEaiBxOS3FKm40RF7jwoUcBJ4NtXnXeVzf94QRinks/40EWDnY8gzlAvqocPkr5zHtB+GFY19wz0NHJ6OenAspzIx
dhupTOk3X/Q/kxRuMyaACC4CnyAETTwf7RIouEdoZpLi19h9pl6LXOC6/Kz7k1UHTrHWP+5sVYQnmlhcjz9MuS9NPlaBdNKdZuED7eHGj8Z4ySeDqWbxMedA4/1lURaZ
1OnYSIZQ+uwIAH5fkRZOQVEN0XFVS7qPH/APwydBTrHzbDgRpfsN9D2w58ad4/uKS7KoMjFEJuVkuZOFtyXktlGi8K+QXQ+b0ucrpT9/ntNWG7mfgYGWd3nuKw1OUxy3
PNyTyt4z3a1t8njGjqxrZ4WBn2xc8l8rxCrRtB25+lZ4IU+NIMx6ywyK2jWU8WysvkUtvdzKTpF22vZis5PCLiUe5TQgdqj9U5E8oAD3aHzCeGlVO/DCgmv9+0YTEOIT
Zuwx39vDciPIv2+YssY9HuVlETj670VAS7qxO38yHm3+k53YAmYcLmeOVFY56VGwkN1PatxQLn6ARD8GGEf79WDnY8gzlAvqocPkr5zHtB9paV28k2kzSWgaChaOzG3M
bPifgW1Zkbei1RhDcOf4FT1kguzPMN9cBhhGj13e9piw7lubAvERByd43dPfb35d9fZScO4rMTW2aOm+sY4Rz9VIEmwQDatSOS6UFBbA5hye2V2TJ/UGnyfU5R60DZkC
PXyMDaEYWZ9qz9uaX47v7DLKDt8H18qzMQ4kaQP292+b+TKlL/GrE5hKbDsjsw1tg2XZS1wGSKlsrP/FdlS0qd7YN+iWSI0zfA+1UPUf1bLzbDgRpfsN9D2w58ad4/uK
E2jAl2KbqYJcHYVkWCpkdggngtzpP/cj9wYG/+HakhaLyr6lAMTJ9WMf+Bi1PTyVQNKnwImUyEZZkTR74W+dl2lpXbyTaTNJaBoKFo7MbcwoOLA6cWdh59L4MfKlOwnZ
xLwhJXN1ZtT6cOzFD87K7qlZ+ZIV8wIb3R1MBfVizlEH7bSZZqbr8C84583+bC7RU4Tz3wkJrmaDiFepi66L92HhgA+/DiM0DPA70xWfkUUFAtntXDDwHHgwesibATUs
VB8e2K9tb3XyNaGbGWJCCVhmezzo/rPb6lSRnp5QpVvtyUsOJD3CS85a7SzIsCE7eCFPjSDMessMito1lPFsrL5FLb3cyk6Rdtr2YrOTwi6a6TdpY8wRG1NQdtunjm9m
mBMyk1zeVfAh/ev0PaMez2O6vTeNsR2iRaEOO3TlB8kyyg7fB9fKszEOJGkD9vdvjWHrNDRxPR/THpXcTSxEsxymhsjLC2SqN3c9bC+k2NbCeGlVO/DCgmv9+0YTEOIT
Zuwx39vDciPIv2+YssY9HuVlETj670VAS7qxO38yHm3Ac8Yc0vCTLNzX2V68A//0KkHTYLZ3eFVgR6Fcq8b8rNOZrTjTXjjj+CPAU9cPFuzbzSdLeFYFkJ07A0w7o0sF
JDUIAcDK/AS2dJ9S0jZEZuvtgYcisHDv1lVcwx9z2M+sYmgC1/rmUd3Gsob+6b2bvkUtvdzKTpF22vZis5PCLjAarG1kTQjK3eqsDSjKOozgD6tcLQvLRAjwnAf7DXtt
yogm0Sa9h4GMq195YwJtiCa8qayw7H1r43fSDmjLEagXI2F/j59yR4t7ltqTMLZBuPCltBUS/S1qyV3VJg10oCFylgIYWfyfnTF4+QxH+jlBLIbatutxP0VgWLgNOgPM
2nFZ5zkC9Z5nGR46t1ow/oQHJq+v4oSY61ZtgxntzmKpYh59ImcWLmj8tZMbSOx81opr7rBw28jEONfnWSRomqPFL+FaUfPZ+60HNcz2UwOTpzLVJ41cmSrdAGazAPLj
VuOw95SQO/1Q7fKPYfQLnGbsMd/bw3IjyL9vmLLGPR7lZRE4+u9FQEu6sTt/Mh5tJBd/KbvpR1MLB1m+WN/eTWn3H9NWKR01H4XUpIQcRJgFAtntXDDwHHgwesibATUs
VB8e2K9tb3XyNaGbGWJCCWSOVxKJis/L9ckaxCX4WCsK41IaCDDFXJQ+j1FRAEcrqVn5khXzAhvdHUwF9WLOUQfttJlmpuvwLzjnzf5sLtGEfU2agFqqKuwROxXQ4oW2
OUHD+DRUQEuLATHwt+sp3k8IqaPKgrArAtAs3nGLFMnWimvusHDbyMQ41+dZJGiao8Uv4VpR89n7rQc1zPZTA/A9H6Kht+k9MpsSKHl/Guw21edd5XN/3hBGKeSz/jQR
YOdjyDOUC+qhw+SvnMe0H2lpXbyTaTNJaBoKFo7MbcybVifS9VKYQawgeCX5h1M/3tg36JZIjTN8D7VQ9R/VsinMbVMrxkDtZnhvClTAtYCShFEPum5NWjpCgqaDqsAB
Rxzn/vuEzVivWN2WPy9lbgm/WgrUKBwzQAydLQ0ZsU2Q3U9q3FAufoBEPwYYR/v1YOdjyDOUC+qhw+SvnMe0H96iX6FHZjwiQ+3+av3hkDfDhHXoLgbC6yQ0Mz+fgjuX
F/7omya14LfPO8Wyvnb/N5DdT2rcUC5+gEQ/BhhH+/XSMSSRfqs1XXNglcLF3fV0yogm0Sa9h4GMq195YwJtiKLhgh/lHE/ZxHkbWDKcIDyShFEPum5NWjpCgqaDqsAB
wFemaqOgW1+yn2xyBKlXVs8ecB+VjDJJGEIUea8W3HdxakMIeJ+UraRTIcOD7H7AOUS31a/6otHwLvNAMxwvIcqIJtEmvYeBjKtfeWMCbYjzbDgRpfsN9D2w58ad4/uK
Eq+98ymBnPzZK0VKvtKblJTI8sPFao9MufaiGUInP/09fIwNoRhZn2rP25pfju/sMsoO3wfXyrMxDiRpA/b3b9DTqv6oACJ02/y2oHBLHtp3NhFJimsRasEAGHoikDVH
L00+VoF00p1m4QPt4caPxvX2UnDuKzE1tmjpvrGOEc/+bX28KY89SEWLT9v3BZPPkyjNbvtloOMTsWlhkUC+Smcde3TX3myCkj9M96UGIEhMdONvhgPnA+3GNhcaQRLn
cjq1mT3EcfitGyxyOtkfuEdsTxHSMe8UaREA9s/I8YFnHXt0195sgpI/TPelBiBITHTjb4YD5wPtxjYXGkES56O9w75b45ssLlK2Ya6nUAMsjH3S+4HJLLna5prva+NA
rGJoAtf65lHdxrKG/um9m75FLb3cyk6Rdtr2YrOTwi7KQ6GZ1CeYIFi4ADbt42keDV/St9Y2RBeMT1cBahGkaMqIJtEmvYeBjKtfeWMCbYgmvKmssOx9a+N30g5oyxGo
z/xqJf/LIzsyILRnCmIBxv98rz9XqKL8vmia1HldUD3iHj0rTxoZ6bRub8ATr+vmZx17dNfebIKSP0z3pQYgSGa5UUUM6KlDTAzAlM78whGUoiIzlBl1elXsVW+2TcKU
OWt/aFcJU3XMQlu7Yg11TNOZrTjTXjjj+CPAU9cPFuwwHaRUJPWBA0rqkzAnZnES4kpNnTsHIOKa8hiutIyBa0tnwuY06IsNIUjRPEV+B9wcu09gZlZiPM0NVkhATLxl
f+9glAybQW7Nv5zLoIcPHeB+8M8gvjijgV3TdA2dzZt7HbhyygLFAHF5eaQuvAzbIXKWAhhZ/J+dMXj5DEf6OajxxpOFukaOun9iT8imrztqU/Q2bk+Yw91eBwss81MQ
u5eeREG+h5Y25UEVu1na4KliHn0iZxYuaPy1kxtI7HzWimvusHDbyMQ41+dZJGia5ASXE3f50sAco+UEGxxv8V33efzMlVhzj3Pyk/BCkJPCeGlVO/DCgmv9+0YTEOIT
ptXwmMx2YQTiiH3kTx1rPt1Y2+MQxCD4kOJNrb5iklJDGzzSOjwe64ghZnKSDFXv+mv3vpgK11DU6/jeiB/lftPtTGHrp8EKdksl7AYphhw4Jhubik7g6x/fOvLOlDM1
wnhpVTvwwoJr/ftGExDiE+/QVPgwlKqQjPX8UbwM8e7dWNvjEMQg+JDiTa2+YpJSxNN+3ZLqeVKEWAnFftNUbMZIlC/HUlo5nMqaWQRjGlYqQdNgtnd4VWBHoVyrxvys
58MdmfxJ/xC/pXizFSAKKm3pyBElbB2DGMBAErJ+S/s3tSbGJyLQPPHNoD8jkrqS49ikr2KDHmwGGOooje69z++qRAUFQx7KLB/ETi3emZb3KJUJrSumrfthvzoHvz6E
hN4LSGBgzYA3AaqvHjYDIx5yDtkxH8HtVPWQw2kMVRMn2XLG6/AEtCF3LozFA0YnZuwx39vDciPIv2+YssY9HgtFffHhvmQ4y1FbQoztc1BHbE8R0jHvFGkRAPbPyPGB
Zx17dNfebIKSP0z3pQYgSCVfT4aV1vJMIWZhAn7E5RgKMwYJnCrjgx/kuU1nY4hlZcrFXxMfhnpVDLIKMAjeXBotccfsdKhpnNnel5ePxadd49uABiJ1jajgXTHnrcas
Nk9/1HF8blZHReiUPVtUGBy7T2BmVmI8zQ1WSEBMvGVv231ERQ/0c1fAffleTiSAWrsnOVbYza18pOFiSn1P2a2WPl3UpB+JWOqJkkljU1dWG7mfgYGWd3nuKw1OUxy3
4lcslu5GOsEdxDClX8x5gJA3Y48PWFiA/1aoDlqUuO7KiCbRJr2HgYyrX3ljAm2IJryprLDsfWvjd9IOaMsRqKPSX10XVnkrlOiWebvy74/SZl6vvVx2bhecBuLOG+xx
L00+VoF00p1m4QPt4caPxqmdNbXB/jg5xgm2NErOYFXfUJXn1TCPRtF9Mzdku29hbBAKYYZoMuVDposw4NVYQ02eQ3dxGzVki22AHXXYq4eXuXc5CDjH1z/6eyKz1AMF
rZY+XdSkH4lY6omSSWNTVzmuBVEyS5AnhRXlrHMUc5iN4j6Ya2JdH4nVrVYys9NhtueDTG02eV391IQuObuPqWwQCmGGaDLlQ6aLMODVWENNnkN3cRs1ZIttgB112KuH
cQcUSummZ3YvPaW/59sRiJF0zGUPIeb7bWQasoaxp06hcaPKGPF+bJhnf4eCu5uFUfFBU3ta5kWZBw0IRpPeIuZc72M2S0iHMbpy7LnrE3w+EVjclhk5GMVNqGoHM7qC
kCcJ0mYVFMDbOgqsQ36yydVjktKNFMTRVTCLTnvlI6jOMywmofQzuM5YrRxCFA22g3+pG+FbCO8oTTvnmsqw61oVWc4yQm3/acB2NHKDKi4b3MtS9qIedjbjdYxCBj/T
8G89ERBHQTzP1Oa9ck3xb0JLXCwojPefKrPTBodWVJRNCJ3arPhhCYVkBWExge7JUfFBU3ta5kWZBw0IRpPeIm1oQ0dQ0RkdyDg6JN3Xo6C5OiQI/fSr6Yjxam9s3Bzg
ZG+WKzR5Guz85pXlIPvKyxvcy1L2oh52NuN1jEIGP9Oy8LFcXMDU488NFnVn6HVwyE2w4FDUgwqXT9t5dt5UJaeb4zBkctBHn0YUz3dv+KhR8UFTe1rmRZkHDQhGk94i
3WGp1YV48LbSwTfm6RauU7eLaJ2f7j7IBdYIP23B/KsYLRKC1B6JVCoDVYvIFLu0CUG5/uvuTyW/jziajhHRyixtyE5kmpdfZAbjScGIrdRyReTbJ2bfO7hxePEB4HhJ
XALlDNNZcVaPyb5pXbwCsupt5fYFgXGhC/j93uCfMHHs7u6BQoy/+7DEoF1ZSbfQckXk2ydm3zu4cXjxAeB4SVwC5QzTWXFWj8m+aV28ArLqbeX2BYFxoQv4/d7gnzBx
44FI0w2yq6YYBW45G267+VoVWc4yQm3/acB2NHKDKi4b3MtS9qIedjbjdYxCBj/TIJGb3/qK6HZEW4o860vxh41czvwU4n3JNGr+5GVWpDa8oItBMD+VqlcKIQoEYAl5
A3YetUVcRYbuOkhPjxRyDEV3M4Fgre/V9WWWD+lpC0c5a39oVwlTdcxCW7tiDXVMHmUPd1ReILbWeeDvan4sJpucyg0Ch0YAGmnQVhu4dkEJzr8LICsgEXo7XZ6gx7H4
R2xPEdIx7xRpEQD2z8jxgXKL4idUk8Wb7R0LCDae1Kxv1lKDHSPAg5M5hYbYvhNuJyuD4VQH9Xondtz4gJL5h62WPl3UpB+JWOqJkkljU1c5rgVRMkuQJ4UV5axzFHOY
jeI+mGtiXR+J1a1WMrPTYQ882xCha1cucXlxCIeW0y2Q3U9q3FAufoBEPwYYR/v1MYpqvrqY7kX3bLozivdzZdLXnLh1ZtRA8i3hs0LZ0cFpnVEQc35ddzJVgSaIaflv
kyjNbvtloOMTsWlhkUC+SnKL4idUk8Wb7R0LCDae1Kxv1lKDHSPAg5M5hYbYvhNu2wh78SpmubMYmIeI8fi6vYTeC0hgYM2ANwGqrx42AyOOXtjqCPTW60nv0frOPqyQ
m5zKDQKHRgAaadBWG7h2QRjTW0XQFxIPisnRbdN6EtW0ouNgomzjPv4xDxjaN1sjJszBeF9yEk5vLXKOlyT+9pucyg0Ch0YAGmnQVhu4dkHLFHBtaCFtSP1ExlM0Pm2J
fxcLnQylypxZnRLmA93hsCbMwXhfchJOby1yjpck/vabnMoNAodGABpp0FYbuHZB+oeKsIRGDA9bK2kB11df3kPv4ssUhKG79U9Kru6tzKC3x1tA77ORJz0JMJAalLXL
wKb2tsycmXx/RRTI0vzGGJl1N/ZSZntrwdbo5o8MlAxoT4BhFhMTECGmG8MrJQmit8dbQO+zkSc9CTCQGpS1y8Cm9rbMnJl8f0UUyNL8xhj+qgFxGwKJKaz7BhKmyTpA
tFED1k4q6Jixr8jUO9Or3WRvlis0eRrs/OaV5SD7yssb3MtS9qIedjbjdYxCBj/Tw04ZNB0m27sv0riZEJG8abHPFjNYkjB26UT4fsKWaiJbYwHhJqINJ6eV0l20N8vx
J8nAK15QmJQUHohwLAlb8FNDHMIheCcpVo90MUXlWrqoNoAioCIuPlGmk8lE3Mh+taT1z16j9AOvLzdPqvvbkbeXO9lYEHsHY/ZLBoUOTsADdh61RVxFhu46SE+PFHIM
9Rcc220qLBp4zlPu0RRUXwlkuKLTfFrQQd0rrvLr4gIjuXNuAhKPXzpdE7SyIUSOXALlDNNZcVaPyb5pXbwCsrLhoGOLpatml9mCgyzNYSOTTkX595seZvqfTqj/rlSG
W0mjlicR8+7GPaf/YWtCMHKL4idUk8Wb7R0LCDae1Kxv1lKDHSPAg5M5hYbYvhNuj+g69/0HrnvS5drhxr3rKko0/2riuczEjF+Nkggdzo/zlKcZNHA1UPtLpFyrgO89
1WOS0o0UxNFVMItOe+UjqEC33DcFlcqpUzxSSseqXDluoGM1YuVBsNSlURnFT0TUyogm0Sa9h4GMq195YwJtiCM3jVZzbd8FqYZsHpA7ebEsEtv8KUDz8TWEb6EKeScN
zpPm025nliyHD78yKnAxofSrSKAzUVCrWouMHcogxbjYIRdMb/ccRPsCSuCwgNkTyogm0Sa9h4GMq195YwJtiCdBPP3F1xfFQAak9KXm1cXDsIlmLsLr4dWNw1B5Cz3M
CyxS2kxcWO91rAKSRBIrhZGI3OU9mrvRiO+NOoP3uLLKhutP56KtseqsBQIPMSVzy4knJA3wljxNNdqpBEfnbWwxtZ5whOv9n/NRwkHoYS67HMoXjBgX9ve/tbOcOUgj
f4cRTw/gWWlw8Zbxv/QIBw2NRPHV493qnnHgFaDNxHHI3QWeJZ2Zg+Pt9myEJVcFcWtLmAS4aXP2xNhwuDlm2sqG60/noq2x6qwFAg8xJXPXqUChQILzhle7AL0urvGW
ZBH5jUfCk8h2i7YqlvL8xdrNPN9cFGk3Ppz+1j52MtgvIAWctCtAOFu9Lf6cmtrSHbJ4AeFdvqGEe12l3g/FHNTwVaiA46lg59pHL8m7XcBHbE8R0jHvFGkRAPbPyPGB
OYChMupP97BfWiV9c2gz8m6MZaZ22Xq/27g0mZ+LpGzswV4yFdfC3u+KIKemjuc2MhkOs+lcmNEABeWuPmc8PLskxEqy4469dei/vxbHcroefTgBRN0eG0u2Ot4Bb6R3
XhGf7mikKVef0telrq/m2psP25WpFEQ1I9FFmobShYBHbE8R0jHvFGkRAPbPyPGBtjpd7zvrRyHcOMEnKgQ0s8wH71xp2I6eRNDSVOhy8XrslpeDdmsA5GPkly2rPnps
LyAFnLQrQDhbvS3+nJra0km0d7dBa2K+n+Gy8LWFKfYIJJLqv2zPTaqFpQ67xstoKFRyCjG0vmqbFWeswnv7ptyTyrsS4Mrz8qThD1+AtO4v5BBlKhL8FipMVMzNsSoX
kgw9fC8RdLWLjRxhZmpsdM+Huxo8izXBkiiknWlI/Eiya/dqnNjWcvNBA70X3G2gh8JeRc3F4Jf2CESdmds6HShUcgoxtL5qmxVnrMJ7+6ZxWBSfMLBx0zMoNbae4BHC
L+QQZSoS/BYqTFTMzbEqF6CNWFICdL2rIpRQR+fpVWfPh7saPIs1wZIopJ1pSPxIasztozThjJhqOhsArxgicNIYntyywk+3rDY+HGOX9MFZJ41Nz4CaHMsRV6/12n0k
iIWrMYUSTqf0cFskWm76El5sn6XPeBngnrXCgyJf0+nCRuDTASprLl6EzW4g8Xg8sKDNhBUtjrZSh02fYLutdTMGs8pcZb1hrWOS8MqzJDeTKM1u+2Wg4xOxaWGRQL5K
+qqS+PNPwrEcVe7zACQJFBAemCj30FWx3/h7eMbbmTKLyr6lAMTJ9WMf+Bi1PTyVQZgtdDqbhxo8EDWCM6U8ugNMe8itzeMt4CL0oSqkaoMF1ExmhHAa8D5yiXQrUMz+
fGy7iQMPYVhW7b9eWXu3tYeVGhLxHI9t81DwOAv5C26ybbSh/nNdB30GWayjQSTOgmcQi538Umj7Pyp7qJU1tLF70n3BsRHmaaeIB1odgNWOjS6WxKBewMIake8VjRHP
RZCAWFOq9vK4Dj/pzfuXgR60Fu1a4T6xbxkNyWRHUD67UX4oSSRspIgSP7/fhIRckyjNbvtloOMTsWlhkUC+ShLwUw6XzVc4mLXw67rCKJ08bwXmiN8+HmXCrxqbA1m9
qcJ7P9ht9EoqVoZqsL19lM1rsKqkhW2JBQj+IOFXQfOjA4flyOWLfuEDU51h/ly9WvSqODQ6YUu4NEtOpojDxrTSy8CUv7GDLrx/7ndWsk5xakMIeJ+UraRTIcOD7H7A
BCzFvS/g/qcYe/Gh9Ji5Ufl10JIFMijTyv0RDoPf4v+giwW5lirtV726Pdzfb0fwkoRRD7puTVo6QoKmg6rAAYtkty6EpijYF5jjKtqV6ldXYHJvzEyG3503fZBpENq5
kN1PatxQLn6ARD8GGEf79cbnoB4hsDmiaIt4bLIfP77/+t/CElmKDXOTNjMWUQLZbaSWBDWDHfTCeJ6DphAmLG6MZaZ22Xq/27g0mZ+LpGz4D2Iig6Wc6l16EzMqT9gx
+RdI6gYv0LEerW55uT7wgPreb8LPaVC2Rt98aooyidp6vlojxiefhl+oiuM3M1m5pmxCVzqEw7JXymLlQNCeVKfR+X1ra/lY1Hh7W0MYaq4ysJ25GTPKWsu5Kgw5yOCn
hG5HWHPey9k6HErrPoCk7NxxdewatfUzEExvqDIMdVNyOROGMSaTqJpudii2q4P2cWpDCHiflK2kUyHDg+x+wGYXctuOlOqfIkVXclPpaEZW47D3lJA7/VDt8o9h9Auc
KCyNXNPOBKDzzPj7FWOnWsBwjoD0TDYG1vORQu4lR5AacLUI4ZtGwp5IAFZWNjxkyobrT+eirbHqrAUCDzElc7bajkcsg+4rA/r8iqRRpkxsGsZqskSgdOYd6V40NmUI
+b59CFjJ7nWtDFD/GHtUhiwuNzcBGuzaaxRiRPWMJF0tzYmOMBL8Dy+Rf8imCddORQjS6Sbpai0L3mHrKh7YWzCJkkV/G0dZ5wCL2HTkyKbLiA9v9xy8Q8bx3UFmvw12
LTP0kdzM35D1SDKjGM0mLQssUtpMXFjvdawCkkQSK4XYgAtLWqA11kZxyorahdZ+Ax7Jf99Seb3JYajTFBdlXfkjTb9kEBHqlRF/xlvBc9v5vn0IWMnuda0MUP8Ye1SG
XrOre/UUPYsUHy1/CBF1nbg8rmjzBv4fgMGzKdjqsI505/LaZeqFaUXG01jNlGLJbz1PLlCxtbvh1BE1wmi3ubGCXg8GZ5B/d2HxMt8MYQoS3tT65m97aQ+k3aqUz048
EnNbunqZum6KjflyWVuem9iAC0taoDXWRnHKitqF1n40UBZFRAeMTv6CU6GqFEuZpoA1NhXCiUdYLgZ9x1q+UUD8Gdq87Ea7cjhac1z94+OjlIywcx6aHTCDafhxrKv9
2EDiErGH25DGUjJRDYcpoQcH6ORD3+T8nqgi4Idg91t6GOWLFq/y44KZtkntEU9UawYxvc4XGSpLOPULaoIGZttOOSKvnlzj+830gy6ICJAEIAdVDFGoQjSgKutiky+d
8KFWU663mkv3H0VnbKJTAU4ee8ibqpy0sEy2QgoEqxZxakMIeJ+UraRTIcOD7H7AP05SlezFLyz05zRTEHRXYGKE95DoyLs2rlV9kpU4USc66kpyaGBvxYMTSqv0ZnT0
bNCAdvpFMR6I5dOZSpmpi8GTRHWJjNVcDCNs8jvzOMre2DfolkiNM3wPtVD1H9WyrV8NP6XakXjvxPYCjOtHb3aVj+pnB4gJ994C5NXXm+u3i2idn+4+yAXWCD9twfyr
DOBwTceL8vbRID9k0tI15HpYEd/45N/u5pUvNZ27iXIEEaDZTtjw21q0vVJhadc9EiRYL6Jh/E8DYKL4wvoyvVG8ALJjXz2FQZ93P8eMAo5kIJ1NRFn/57Sox3JK6jFN
BBGg2U7Y8NtatL1SYWnXPRIkWC+iYfxPA2Ci+ML6Mr1RvACyY189hUGfdz/HjAKOnWhAF2eRc3poa4ITM20wdnPrbEDm6GZP4yo0u0FxxN6zGcoZu5YtxJlU5cQhl9FR
/FT73LmvVVNoucz2CoousbJgiPFF56jEYZnzgKBiOCma89Z6nZw7hafcxsI+qCS4bNCAdvpFMR6I5dOZSpmpiwsvgHCiz0SoFamZ16/LphoFcetbs6j8neFFPqydZH00
EiRYL6Jh/E8DYKL4wvoyvVG8ALJjXz2FQZ93P8eMAo4yPU8GfdaZZ8KjvDOwXJmX2lbPfqvRFH64mQbwxBOPLaUZ6wW2FvHMGzYOwXv+GRd5kuGBPqMBzvcw2WJkFXOA
cb18/uFIkTgCAM9tsGXXOEWK9Ow7f8eieCONcCmTQFvdKvSRnYvPVX8TOibl+OscWTA2rAsQvBT1MFPb0CpP8/G+YETwrBdrNmLQ24ltmEf+1tjDCM8z9+66f72n7sLz
5vCdy6CQtYl3Lh3iVpaCXnVQDzBFKbLcrhJuoD6Yjnt+/OjPKb2IhLBGlz2LQSh2nZjeat1EMVfEYMQWbyk+K7g8iQBKJ3IjPqdN7OX9rG3oXkZmqZxds+z3xmT0ywVZ
nsoty9cp7CMuTh+3wJJ14sqjOJ1IHNdr2ulltZdPu58KuD3sOLU7bVtHch3yQSKGjeuO3O1+yFsRCkprTyZfaxxHg5D2sVT64/nIsn1dOReoUsotFmZbA66TZxWX+JF1
hN4LSGBgzYA3AaqvHjYDI7v5LBZW/9SE6ys4MbKm2Q0R+YWp9P37wXyrZcqIMPcPAxvyA9bgNQYIbsX2j0snuYvKvqUAxMn1Yx/4GLU9PJU/TlKV7MUvLPTnNFMQdFdg
7aVObc7o04onA4Qns1mM07hkBIWjG6RweLyLIx6mV+QLLFLaTFxY73WsApJEEiuFg4UrRYiGO77dRrqhbNh2Rt7YN+iWSI0zfA+1UPUf1bJOArcph+mLWBke1oIiMnap
49ikr2KDHmwGGOooje69z/MOHrefbuYXqD+n9CuCHf4XXMiFnRoBWB4VkmhT4TU8v2B3hWvETFu5jWuuoady3ljlrTtLb+N4fsBGPobszps21edd5XN/3hBGKeSz/jQR
jt6/YxTszPZnwBicSafn07eLaJ2f7j7IBdYIP23B/Ks0AyDydX611xjP3VcA+E2w3W7CXfAnjRNyYoElAvGip09+L3KtJukqBcliLCbmU3/agnAn54NtcLLArsZhghW5
7OwXagq6jpxtqQJgPOfoTibuQRBxrPHb6a92ceabR9cqQdNgtnd4VWBHoVyrxvys7FQpJztEMEN8/pd1b5bfkEdsTxHSMe8UaREA9s/I8YHB74hcOSi3GuTL/y5SpJo/
yogm0Sa9h4GMq195YwJtiC0IR/qz9CVDIaHhbtvCp2CShFEPum5NWjpCgqaDqsABNm+PdWXSFKFIw32EVhUSZ6mp1moLM03ufhyp46yLNKtDG8FYtsToNw+ZZH2gkWrc
yJ2lI5RVftkwdnAnvz7XlIydP6XR6e4612NIproFIsJJYySJWlq+qXWZJR8Pwqb0VkoRC48RMHqbCN/BQB51GMqIJtEmvYeBjKtfeWMCbYgvzCMMZTKt5zEGzRWF/guc
49ikr2KDHmwGGOooje69z+4GEY0AZsQmiDkLh5sdTTDN2zbtICS7LPpyY3GIS8JXyERaGp2S2i2zA46pdBcLQcabgt3Uh1uFDtAxGs5UuqSQ3U9q3FAufoBEPwYYR/v1
rQYFqbYuSdkIIYozOjk/ZW3pyBElbB2DGMBAErJ+S/tXQiPwQTBUGi9dxE7ltOFbzAfvXGnYjp5E0NJU6HLxem/yBEB06P8DzXscE8wFd/LEb7O1r0cxPqEjb/MHm6Jd
rfY8PN61rfh1p2aHfrG++ORQAthhvjwfTu0GwGsunFUqQdNgtnd4VWBHoVyrxvysRyza6YFfeG2stSyagNfbdBhA9MAjq6BWRvdSWqU6Uhyp2ablVBOS37XWbdGSh7V3
J9lyxuvwBLQhdy6MxQNGJx6qJqlfMQHYsMFjbV72eI1fHzzWDDhjeiTAHtl0796VRW4NOniqJJCvdbitsYK6i/ejenr5XTsagrBVvcOvbYvI1B4Rl4XeelI+3QHBR4xl
VuK8O1Pioh0nu15svwe8Q+PYpK9igx5sBhjqKI3uvc9lth1YPbXvQFnuMkx/Jh80LOVaHV6j8IGu1J9SAxTFpvriQscXDVm8bgAFhHJp2wF1VmNgm6BTwYg3q9CWSMKs
rScydRfi2swJNgabVvp34FXjyubL3fuBWKgCbq7S1AXCeGlVO/DCgmv9+0YTEOITUBu/BoqljwxSurHe/jCAeIISkwivqSoYnUOrgX1IMwdFwigq4S8Q7Zrvm5RchTdk
+RdI6gYv0LEerW55uT7wgIAdaUYtmNnhnT3kuJODdSHGogtdCHIGbGrP5IPM66x8K3jLMlHAzBu0+n689gXkETltCLfeHVcvT46kOw0APMvxjPpa23CBSu8nEHWbkDh9
pz7D2U0EfKaDJX7azPYh5VZ8WfAVO88MQ3+vvJ+o8+945GrN/zKCHnQRmegt/TjakjoGSculgxdn5ceragj3J69BQR94XczNQD4KancGBk0yjgxVQRdF2SYoFghbH0H5
R4mNi2v1fOFVtotSrTdd/FvP8r7aNnJR79ZcXZmKa7V+HbtE5dcb4p2jdJZV+0d+LCHnqKPu/nDLVxcYGsyvULeLaJ2f7j7IBdYIP23B/Kt+i5pXc03iDNZ9MuId5svb
ITnqnAra0AOO4jMQqxAZp2u+C8ttpo7qFoCvCK7csmjckujMgPhT2rxvYW7pJj4vqqQzFdZph0IpD8J42MVM2IqIYpTewKzeLplZfK1UfUU2/biYwwwkDGpP2ocV3bmg
UaLwr5BdD5vS5yulP3+e01M1Bd9kTFX4KLQCdg0x23ciWeljkw4RRBljmPbnVg4QlltXmzjdkXVvf22BQHxrKIC3w6Vje4bzzgcn0rApeYdRovCvkF0Pm9LnK6U/f57T
UzUF32RMVfgotAJ2DTHbdzaMISthTtrlwI8Zsnof+OaWW1ebON2RdW9/bYFAfGsoq9Hi3CJZpkuTeHKnxsT7q1Gi8K+QXQ+b0ucrpT9/ntNTNQXfZExV+Ci0AnYNMdt3
QXtV5CULKMauCgQE2V5YDJZbV5s43ZF1b39tgUB8ayhAOK7KF7adhwJDQlqUGZazUaLwr5BdD5vS5yulP3+e0zf7nLqzGFxqMWvJtqcyBP4lS/ohHHir/d0TIIgLDvxv
cIkmLY/wBi2vpI9gDYHW2Nm+PHV/FbC90tIIxYiKNoG9Y/9WeXmsZvBwBcXrxmapowOH5cjli37hA1OdYf5cvZXWxDShVgEo4zV3lq3Rnw0OKCjxmKIVdLpm+3QLvv+o
jc2y4T2uCHOtYYwbg89ncIHpNTsO8V7skdivCxmxRIlxQVnaDR5XaZ4sfQI3j500cUFZ2g0eV2meLH0CN4+dNHFBWdoNHldpnix9AjePnTQhPRrlR+ySn/OdXHpm3UHZ
rnJTJVkKdQgNXttzOfJ/7LZLkRpOXwNdvUQbhAeIqNQM4yqFlwd1fLcBIYIgC3epcUFZ2g0eV2meLH0CN4+dNHFBWdoNHldpnix9AjePnTRxQVnaDR5XaZ4sfQI3j500
FDm0UlsBhCZQN0GGwKwvYq2WPl3UpB+JWOqJkkljU1fqgyx5D6+evNVTyCHKVSAX3tg36JZIjTN8D7VQ9R/VshTT/s5m1XIByYdpgKEBsK/j2KSvYoMebAYY6iiN7r3P
GTnO0QFtsE3+ylFrlEFnAFWb1AVjPSEku9JU+oEDnMS4fSv+ya99oL0cNfNbTLQWYbpnK89sEuQHsV2lKPTy+uXjtPz5HqnHIwXEcFgwR2/iHj0rTxoZ6bRub8ATr+vm
YOSsabpsQaU2VV+VGBcfOdUpl1udsdK8QGuruoiHmLug6cujBu84EncAPKip38q1wASIya+ayT6B18GbxLUQhZZbV5s43ZF1b39tgUB8ayiLVmyZ3vtpWhaq8rkTIF+5
4FYJm/PqkaapdPuFv4moVRk4bU8CZJcF1Bon/sOudFFRovCvkF0Pm9LnK6U/f57TsEwZ8i7OprjDv+1oU/WMzEuH+/v+3XW3eShF/6MxtsyWWeyuztfvCdReXG+sovXl
fsOBwQh7K47qdDLz4Lyg4pMDY1SdeLiPAfwqe+HuMMDzwz2HAViKzVNc/IB3k4uDa87toigUy5ivCQM/ptx+krTgtmMTPgqj3kafkNwo2HzLhjq/aSEOgZwfPiTu+YD/
VZvUBWM9ISS70lT6gQOcxLh9K/7Jr32gvRw181tMtBZhumcrz2wS5AexXaUo9PL6i3v3iJdIswaQS1321OYx+xjAAbDnCR8KX6quSKwIX3k712WCVXDEUzcr3vJN/M3r
g7V/SY3UW2i0hYydn43bVaXl0UNAFO0yZl7MyFhHAJHbTYH8SiMpLaYPHT4HnXSsUaLwr5BdD5vS5yulP3+e07BMGfIuzqa4w7/taFP1jMxLh/v7/t11t3koRf+jMbbM
ywoYj57aDZL7xNpDLJ0FmzR/bYSs7JlG5BokmzEsxkgiGP8sbF0njmT7/2yI8rkqYOSsabpsQaU2VV+VGBcfOdUpl1udsdK8QGuruoiHmLuPk0mWtkbi1W4HOoq2Jv3M
rn78wZHKVIsCS4UzZcMAZ5N/fz2cqgMRXVPkQ38/Wj6uhYu61msoBRfZlualkmykDwRuDyzPXdDwNDCYf1wFiwYeADa7GPxP5A2lQOZQZoYg4bhbVoVNR8l5+tmh9qcW
sEwZ8i7OprjDv+1oU/WMzEuH+/v+3XW3eShF/6MxtsxMAvq+RjJ4hhZsIG7/CQi3r6uswtH+RPHhIjhnu1vw3ezzOnG81fWaUX2+9m5kxvemvS1HN3NmjK52oHu08mB0
VLtOBSFPTuSVSuWE53RV4jZzn3b0SH4lmCEeueGMngmVjoUfYTp0TiaZk3zr7jDARMe0g7shdEuSAHNcBohXCRfIoaZGAkH+NWa8lzShduKShFEPum5NWjpCgqaDqsAB
yPJVrGexs+hGNBnPHZnYSFN7Y2qYm5mE9wDJq7eb9duEyjZDhti0G7QIyeyoDMxJIUj20Fdxg5KMSTkjetcNp6fSm6k0oleo07JP8BifKH+7O48FOALxndLiPIeJrurD
JvW2tSuSh49MgIVy8e14N3ZQKrKRyBb9Un6xJrR0waYuQ+/weGHIlAJI3B3Srnkpwyhknf3OC8em1KN4gx4MdBXhYKEk1w4ZYCWc/luIR0mBxP+BwMsHPKxhxLbF1Wg1
J+7uG/2jzz4B44UW+UrOn8J4aVU78MKCa/37RhMQ4hPggxNFlR5Fj0oydnAJ+/qdPDqzRMA3TXLmw/DblS10MMqIJtEmvYeBjKtfeWMCbYgea9a94O//9H+vzG1nuWA4
A2tMMHYE6/PWCXFcu8kowkRpJBMRuyVqdznXv3ai9WdrvgvLbaaO6haArwiu3LJox/n/BKQot1yakwsRSipgn33cwEIMC2WUH+Rh/GllvStLZ8LmNOiLDSFI0TxFfgfc
gcT/gcDLBzysYcS2xdVoNTi32qU1ndRNgYUKhXASl0ocpN/f+378VAmYXpJwDf9SkN1PatxQLn6ARD8GGEf79aeHS1glvnknBJ3TO4lVPrENg+kNNc5dAh0+Kmc5ztqi
I4vtb7teD3cMqKyC/5xtfGu+C8ttpo7qFoCvCK7csmjH+f8EpCi3XJqTCxFKKmCfPvxBUgCXdtYWr9vqq4wv3UdsTxHSMe8UaREA9s/I8YGk5MnZjnxwDkv7h7Rj70GX
ecYHIXd39k3jckq5ea4jps1rsKqkhW2JBQj+IOFXQfPiHj0rTxoZ6bRub8ATr+vmCb8jfIKDgB/N82y9DzCQG48voa4gfNiepx8vlZOgq8yFQHGixm8RgSZyxe3oTWPd
ZdVxo76EJm9C2itQjolVeHKB/2ChPrHoy/ZXH3DkM1J1zbK3YLPpMnJ4CEyJoDVPw2JwE1+YZvUiXkLJMKSX4PGWV8c1Z4dymM1VB4TSdA0AXyX0MWJrztWtLn3j7LcX
2fVFfd70gPzQ5dZ7NDfaMPRk7VT0y6Ycs/C4OHtGB0dfYzzkrDM3HkNXFCxOHDPN4FnI3N6XN4sRjRu34PN1nymO/G8ONsRIAQfXY3ibsLYOPxfDZme2xphGob9s2j7q
saA+QPhvOAzum0iLzvYspKZsQlc6hMOyV8pi5UDQnlTXlQDEfOuzT8oVErYyLm5OgUHmPA7g56a4ObVTBkW9kjlrf2hXCVN1zEJbu2INdUzfoSDrLK8yDPnm/BqyjG0s
pLQ8TjYxWYEoIPaM5TM9K4wUpTZZQPnTiEM2ojsCEBEpjvxvDjbESAEH12N4m7C2+Ufxjg0bsA5wD+uXfKbmfuTr+6U+JPNCp6/679SUG7SLyr6lAMTJ9WMf+Bi1PTyV
iI2lGGkK/dhasys/iD3Lm9IenNeLWRUe+1SnaMuooBuQ3U9q3FAufoBEPwYYR/v17UBMsqVRg1xEIh4albaQKX0Lzll6Waf0QLoMH9x5jsR1PO4SZ+ZcUXYQ/ySlbkmo
bBrGarJEoHTmHeleNDZlCKoAc6zXMoCe0JU0SCFrArX5G2XXEocUmNbAoVAO7JFvrZY+XdSkH4lY6omSSWNTV6ZsFCKcBMr4hUTUkshuqusZhFG4YQNBJst3y2fMjypo
BXHrW7Oo/J3hRT6snWR9NB4+8zBVmIPbYuBTk0mYmab2UkrbfmSv3FVAZh9XaQ5Sl5DxT7WlChXbI9ZMd8y8ddP4miryGw1RNFRbRbhuawD5ikFOhGAKKFpRVlGU1+2Z
X9i8LsBkEZtJ/XQElOz2q8qG60/noq2x6qwFAg8xJXPU/msTv1u6SwE9Zpcmy59iiIs66ZCDiM3Wal55Z+PgtOqEXCsBgq2TA0YDRx/RJHgw2A6OEX/MFUVLSiPqrUI6
XHi44zK3yv3MziE18IUjb+IePStPGhnptG5vwBOv6+ZpeVXWLLkPMZTtE6ZLXZaQTM1e/GU6ZiEDmfUq3OvCcrT2N+DChuuYPncSOz5xuL/s+jVMws7Ne5yQwh9O2Q7l
Vdf/k32siq2iu2NUSA5CjFOVXXPgGXpcJMw1T8ZqMc8yNSLjnNORA2yWw1gaj7ayNtXnXeVzf94QRinks/40EZShnBkvLCnBjPn8cDUhyCO0NmGP37v5Nd9f5TgXgvBz
X3pynP15kpxKrmY6UizunV3+SSQ9kqGj2xzK8MLr3hg21edd5XN/3hBGKeSz/jQRlKGcGS8sKcGM+fxwNSHII0oaqQU9QIo6ofRzHOPl6wHKiCbRJr2HgYyrX3ljAm2I
D/JB6V0a35+swecoZZfjo+NyGKSLWlN4DJWJ5QIkJ917ZgjxZztcI0kcczrv/GD85exER6/DalZg/SuC4jYOSsSzjFGG9WIEclybeO2ZHGIhxRWOMbRrgLEFqG+wx2CD
qI/IhTmIrnL6N+rCwoPtuiA/bgm8v/rw3kYbia+lbnz68PUeBF4WzG76U96jna13NtXnXeVzf94QRinks/40EZShnBkvLCnBjPn8cDUhyCOSlZw9sszMwW6R1T3SSNgR
xkkfUWljnq63VgXQAwYElyHN457v+YWrapG5f66+ZOiNavikZvNew6Y8R2Sok/56yobrT+eirbHqrAUCDzElc/g/wrMA5XGEFGMERCl+4AeK02Pn73xnwpllm91h70ub
SZSALGlZg9ttmz7R/BtS3f868AlTV5FyP7uSAn8i0cfGSR9RaWOerrdWBdADBgSXIc3jnu/5hatqkbl/rr5k6JCoLQuqG3EFLEy9K39sSt/I7XRiUaobfEspOor+mLHf
0/iaKvIbDVE0VFtFuG5rAJEQZXIc4H6GzlckCSqm98QeL9smrGapvMMlfTHHZdQyVSfznKDSXN9/6wGFgAvGLDdjVJXihNkWIFjyAAcNx20FrHgZXGWY5g3Kqp0jfXYp
+XXQkgUyKNPK/REOg9/i/1osW3UCXQQk3RlLOknwdd1Zfu6xCAv67rYOW+qIlk3NEAaRPMwj/GUniX9Y96PGwKd0Lst5mm81N+MYfvzWIObOd6lEFhb2jGDc2BmFtg7z
rEHexARfYqFL2KVM5G8JVEjyO6wFpfx6kbNsb93UVmtvf+NaBIJkC4UO8SJcWxdjvNbMIWpYDe0onZyFggiLUTbV513lc3/eEEYp5LP+NBHyBwCwFKqqhMxUO80gmGxS
GTRWlTJHuSNtvjqjD0OVn8ffiQgw/+Yu5/uIb/iBxMw9FMJguPrOTK8Rc2O/d53PJX8ANqHSQ8N9eUIUjNmVUTyHltK2hvepmExZcDzyGVe3i2idn+4+yAXWCD9twfyr
Xq6y7r8ZAAAowKM0uWS1OWLizYXSBW7kE12IyRQ30TnmtrhU5L8tJIWu3vlHxNo9gnDkM2W0BCK2/GSLcRfLJZ77H1bOY5BBVkIV783x11K0B7Bmw174pKxn7z5QsS8z
1tlTSSdghXQdbNDWXjT6oIz++dRTErPjK3GLYFlEFJMTL35kR2ttW6HfKDfJF6mrRQeZghvvbzto2QWmwvOUnYz++dRTErPjK3GLYFlEFJO9+iIhGfe3ct4hZ2mAhhNM
lYzI1XYLJ45Nv1Uu1tMB94hujoyFqHwUKq6iIwpEH7JvYvGKctXO39J+WzGUcP621BaDY02xSc5UF/N2FRiJv1Gi8K+QXQ+b0ucrpT9/ntN+a9U1LPJ1dY3HilVwiKnS
AsxeiQkM4f66WpvA1Pbqdn+dYoI/sZiZrQOkxaClG2nKiCbRJr2HgYyrX3ljAm2IWixbdQJdBCTdGUs6SfB13VEfqU9BaYtVyGZBEIWbagCtRGGV+QtUJLhmsA/vaXzZ
yogm0Sa9h4GMq195YwJtiFosW3UCXQQk3RlLOknwdd3TVmRz5h2ONhoOQv8vSWS4c2pLvrC9BGP4pILNsvl/u8qIJtEmvYeBjKtfeWMCbYj4P8KzAOVxhBRjBEQpfuAH
K7LDvbDCgWLJ4dompIXXMJmh1xl3yL9PDeSpUkcYeczcD8/GBBhaBgkLK12fVWpRlzBX5I62oCKZJ2Mk+Gl+s+oDQCbGUkBZXVnjCrlkvPfKiCbRJr2HgYyrX3ljAm2I
+D/CswDlcYQUYwREKX7gB/1MlwPwec6MH+VIRqp2C57KiCbRJr2HgYyrX3ljAm2Ijf1/S1xKGEgusIC8ZJR0ZTICLXFoGdSwulyDD//XrZdRovCvkF0Pm9LnK6U/f57T
0zxcTo8fEbtcGyjeqzEBM0oJhBXvLAMf8iIrF7MGwL8lPo/ncQbZve4jEQzhnKmzZcFZF4eX9X4du650aJrWvCiVtZa2pZC8ooY9AOPn6Eq2lNeSH+3TzOT1l9K3H/50
dlAqspHIFv1SfrEmtHTBphBBoc2ZztDDOfCwfqo4NSqQs7rpXpCuXaOMheBUUBbLJpz6cFFmfbZq5nb9+T7P/t5vGkerRUlChsrGm3g97sY66LGAj8uziOICfdhxX2PH
4BTcCD8LSOsXr9tM0SGgLHpBdfRN5/hMUv563Dt7aWmWL8U3VOcvBVIKavZR6GyZ9J+7dTm0QUmaeVVZG7nKW8qIJtEmvYeBjKtfeWMCbYhaLFt1Al0EJN0ZSzpJ8HXd
jyFAFcG1iVwv9yIJnu+RFfEzCcJLAM51HsKOUktLISOWL8U3VOcvBVIKavZR6GyZFyvdwN9Sn0T4jVB5ir3/RBudMUpOvEviX+pDvNsbFklvf+NaBIJkC4UO8SJcWxdj
FyvdwN9Sn0T4jVB5ir3/RD0UwmC4+s5MrxFzY793nc9Dl2PUnmVD6WlF8WqNq5oiizIGTNLnY5q7QqJWzp3kSCmO/G8ONsRIAQfXY3ibsLbiGbs2iE8vp0Vh6D7g4pBg
2Rn8+lPCXvmGUo9ONE6WpAcypABRL5m9FkWTg8sx/bojrWuO/qdiISHDbRC8MJz85n2BnGlJA5tub+QncYPht0UHmYIb7287aNkFpsLzlJ2M/vnUUxKz4ytxi2BZRBST
Pl1ln4mX0UDelE/1pUI5mJ5c0Ft69dfkWgfh8y5E1Ax0vqLrMYA3GxD6ZC+Z+5alcEck5tvboZNKlU39STEJHjlrf2hXCVN1zEJbu2INdUytzwnkvjpM6GtxpFos4rSg
5CTQDqspM8LCxuOXnkX+5e9QRXlbAOythLHbWs3xco3TPFxOjx8Ru1wbKN6rMQEz+BoFo3ztFlX7o9QR6QjBXO9QRXlbAOythLHbWs3xco1ZaSdDACS5FUiRb927QIXM
jUzmjB26sDLEPx/WDcn0AO9QRXlbAOythLHbWs3xco1+a9U1LPJ1dY3HilVwiKnS+idW6A6QYeDjviaI2VOM28ZJH1FpY56ut1YF0AMGBJchzeOe7/mFq2qRuX+uvmTo
ylyTNP6rnSaCnKtoWj5kQ/l10JIFMijTyv0RDoPf4v9aLFt1Al0EJN0ZSzpJ8HXdUhZ0M+SsZize3PSfynJ2JWXBWReHl/V+HbuudGia1rwolbWWtqWQvKKGPQDj5+hK
jkPC+N9p6iZ4nHmgs+wcsaMDh+XI5Yt+4QNTnWH+XL10vqLrMYA3GxD6ZC+Z+5al9Hinjynk20bN17/xzgMPFo3r3bzM7n2Lz04uEcMWtTKXMFfkjragIpknYyT4aX6z
SPtckLylXInOvayMasQMau1+Sa0ZXl/IfXIAa9wXwFHzJkcEQa90TbDj0fzy3HAKfzicU30/6Hs156zdIwzOQZBQwp8iygKZH8qQPJpl7vDtfkmtGV5fyH1yAGvcF8BR
FBLzulbNQKP7JIqbTUY7hQjujVh2gxpAKN0ZVUoDxcviHj0rTxoZ6bRub8ATr+vmdL6i6zGANxsQ+mQvmfuWpchMmCqSqV4QTQHGmaVt9biS3aVzLPlO/yh/9eGluSjB
vW8bCb0YY/2VofyvieOuBUbdcqu/09eph2KdoVQL57QW1mNzSN5+r5TlVyURsSBCwFCo/m34ZiuuKR8NoetrarTKkTNoFF8+Qi7bclRAeJilYtSVSeprOjrNEHarp4jU
dlAqspHIFv1SfrEmtHTBpiBe2FY3gZJ9AMRTI2JA3ZIwsaK+RPg+t/howUaVP69twmjntsn20ecoemcNsCZ0v/l10JIFMijTyv0RDoPf4v86m+gYBqbWB+FIpSLP95ut
xiGZOJG7bk1MwD2rntdQFbuRGy5TzYOcT1z4syYYNUWzlBq9zWR4XHyL8Ubt7MAkYyRqI+xGy1b0Wr3qR4vhkjkko8HdCdrJOIhYZmBqnXFeDdUyu0psgZiVKRwhJSTG
p3Quy3mabzU34xh+/NYg5kENpqnl/O4fqHNkD///QoSc2YkUvAb9dIgtxP90vDF4l+mdgiy7utQBqQqRxXMmHaTdRwJ5Tx8WFJMO0NjePDSumldEg8j5Na8B0W+B7dz0
6SFHYg7Obz2p/PumSAtYiUTjc4Zh43+1knPWja37a45bMbvTHjAYuulxkqblu0hcn4F0wurjdYp7Lpc6vV3dp5R48jfl0YpeL9ojaEDo/DrWAtqDMcZYJ1v3wvbnEAXD
Mp8/W3lp6icrdpU4NrI8JiyLp8dlEjQaBt83dbKwBtXfNAcLHl/9LLsEFVWZS4gTvV2RLlIT0dMefPrWUrG8UdnrWg5RxtuZluTv9obzuma3i2idn+4+yAXWCD9twfyr
Xq6y7r8ZAAAowKM0uWS1OfBR1BZNKhz6FdYesVJpp6CjA4flyOWLfuEDU51h/ly9Ye9YKwduGZrQiyfzHq8vUe+NYLheKLn7290oxDGDjcqpbR5u06j8IwpQL+2x9m0z
foZjCXBvfNzrr/+7oX07KEMpmpxCy+LVgZlIpneFw2kWd75tqLe6NHEQsFSWZfL/qMe2b8PhvEUlt7ku6UKISlGi8K+QXQ+b0ucrpT9/ntOmbBQinATK+IVE1JLIbqrr
pW0sJfcwwYzSvZr6uVpjd1Gi8K+QXQ+b0ucrpT9/ntOmbBQinATK+IVE1JLIbqrrVy0EvLwFt5w4sfet/MFRmOIePStPGhnptG5vwBOv6+YHSTmjO/cDNyJPckQpInZP
KL2sOf4VITDO7C4JnQPmhLeLaJ2f7j7IBdYIP23B/Ks3hssPm/UFPYwV+E4CIWrojy1fNpAI1fTR1+Upb/cXdsqIJtEmvYeBjKtfeWMCbYgw2A6OEX/MFUVLSiPqrUI6
cO3NbkQFo7pnxLBEaafpdcqIJtEmvYeBjKtfeWMCbYjU/msTv1u6SwE9Zpcmy59ibab5KTBihs5iw8OI8NDiyvEzCcJLAM51HsKOUktLISM203gHGKD32JXG4q0CvP3w
lfxyH1vNPX8uh6+NTBiNJWMaMEVH1Tvlq4Mn9KQKHKVp15WsYQ+SRDSbr72w98jZoGaJUP7G8YKABihfmmvNrxSDk3t+Jcqg+Ja7T78RX0v5GUGjtZIu3hHOSSK3Mbqj
Zj+Xk0xmYkm9HtzfsRCr0SY2IBIoofsWECJJ+aBnw1X9wpyXHXy7BUCgJK4ObSteyN0FniWdmYPj7fZshCVXBaj3/NCfBqFNP6QRIurFFbX5ddCSBTIo08r9EQ6D3+L/
Om3fQ4i3T+D3CFBGpHhL6epDJGdy6uREadhz8T828azd2ABwBFoMt/aG1eYjCq5yZwD3BkmqSV+SdLDSH/Px+A0l16k4YALBOoewP5d62X3KwxYvfqeZCFI7hdfm+3qK
jPry3lrPEy6GKRGe1Mpz5KcSj/4XWo523coRqaaNw0SH9Lm88DJQ7RASk4D5tjacv/FGqm51GLcIdQ+0L4nxHwT0+S5To9oRarDGytJCsHHo/vPFI7zTx1My4M5NA34a
XCi7NK8tSOz7JiiFqGTHTKOQSdrnhrJxLP8w7bomDy/pkc7wGx/Sr24yBuXN3VNglpOh2i7aSVMN1UQ1IJ/l8HxBEWfo//onubEX7O3Ur9kTGBsPh0+xyGC9pDQ5Q1k/
ZMo2Xqu7GKY96SWjjaDuDubjrWi1ypMr+hPplT9aUBnPPix9ExUWb05b+sTYp+H8A0Qa2Yy7ZvpDLkamXwz7WTc/8xM4vIXLdH2oWygd/EYqPIpy/61JjIH00Ma5Ex+j
Vw6q5wxBoZTq+qMtUS2M3fUJ42ZvbyXjaDfltAmQdThMnyvBPxs/AhZBImEMSdF3o3VCYmmijHcV6tUzaYjEdt4fNo1vcPRazMfPiXIJcFTxxueGY24W74fnS7qW0LN0
sxEouxCdukVbKvdhNI1hC9K9VN/mYtbtD0GTb3ykcW7Shat1UtxmpKKXko4Xg8nYwNsMgOqTz+4XKK7j8r7aukHgLa2NWwmv1/FExJixFKJCGsVGQYC/wbQH19N5iRSk
lpOh2i7aSVMN1UQ1IJ/l8JkAr3aEzsMGvMMdO4K+pPwVy0gpRnyWfOnJkf0UDJRwksdf4S2289LuxME3tMxVSll9AXDJg5vGu//rgcMn902jkEna54aycSz/MO26Jg8v
MdK987FhFR7dbMhMth6B2nSIYxKkbZw9mbeMJaGd8xkGBuwdXD+3FIe6dJd+qOunIhBnNa0zLVwUI7TAYFYWCgj6besWU7X5QfINhxskpga4Ez7eSoZc7vw0ZIDzp/fH
YT6T1RYoiuHiaFGFkjQh89YtUBuNOg3xYtePaN/bCeeH9Lm88DJQ7RASk4D5tjacoLNpSQe125amuK9KAj83Q0HgLa2NWwmv1/FExJixFKL7GlWVwHvOqxVq/O5a07wG
lpOh2i7aSVMN1UQ1IJ/l8NhZIppfGSqqn3VFSAm/SgFB4C2tjVsJr9fxRMSYsRSiNx5hlND3O4SeMf3wfUNL1ETViyAvwRB0UOJhQP8TFyRhPpgEAvbwQquaVd2OSwks
o5BJ2ueGsnEs/zDtuiYPL/YW+vo8xeKTLHCiySwIPCWzESi7EJ26RVsq92E0jWEL95LyKTM5sCSWJnG90wTobEHgLa2NWwmv1/FExJixFKLrmd2j4wTzEok1VcN4VKKF
ek/uFlWO6ekL7VDHAgzZ1+j6I/nPT6nY5WrxW+FDBb5B4C2tjVsJr9fxRMSYsRSivRwNjpw8zoAp11FLzGQ/rsP7aEJjY9mNdTs1OE+ZrwYI2w4e/Ey9NsLeiHgEGj1q
Xd0Ta2CgosxZphIEyCfjssss4xX8LpMhpX8/fpzZslxhXZYCnYUzYF9dsEYYCXexRzBGq0o0BAuBTbgYRWvrZ12ltwWj3YUXwxdykGH3WhwQewlkhqQbxewt8bD5VB2O
zQhme1rVT51YAjQhc34iHPyu6N8NTGcoy8BoVdqYBEis0t+L60wrU19YVzNUhq/+divg9s2mij6IKFVIuu52rBMnlw4d9NFsiczd56Y8LO7HsuOo3BMFAWik+9g8MAFy
QeAtrY1bCa/X8UTEmLEUosLEoobQprEtc1fi2ElRdy2Wk6HaLtpJUw3VRDUgn+XwVoDGQ4Z5/4G17gKLkJoiGEfWoFdnjMZ3nH2WCYsv3RJm8ax/ntJyceCO6vrQp803
I47yvhpENBhsJ/mzRDvrbkt8QPCFuRaOKH8veCt/T6NkCyp5D7/RjJ4suPrnB+MDTCz7sFRpMKaJMLB6MZg2WVwzE5dAZtxPTbATG4pKtPsCPb8bINWVrHhny9e6fq1A
qDFcCMglbVIixlKe1qzSjTNvbxXnG3L1F28QeAuN8m2sI406Fybs3/N3t6u9eQjnE6RvJZ3r05z2iXufFyvGhZmLcZg7SL5N+7wp5DZwfBW2RDBbAvrLmgC5R6ziboHe
JUR5ntfRpatTQI0uo0GV9KzS34vrTCtTX1hXM1SGr/48M+ERnW02j5LnfogfDR11OYxPzTbGPIn9LjTnTgyo1BJYgstdnSXBRbe506+7JeRWRAIWpqPVBaSoW2sIr5Y3
KjyKcv+tSYyB9NDGuRMfo/y3g/CmeJUfzY17ZRZuwtC3Mpz35qVhnRXmT2qnELXCh/S5vPAyUO0QEpOA+bY2nDLbQBmY/suCMfKeudfTVstRB+ZWjNKYkGtGUAR9EPkM
LUP5CLm5KNGqeVDs0BalFCe9W2p41KOXJ67Md8oc0eeHlML2byA5lg5y325q6VIZf7uq0+dYLdYoWzlPy1DDXx8p3Wm6VgmyKim1rxI542N6T+4WVY7p6QvtUMcCDNnX
WixbdQJdBCTdGUs6SfB13XVDlE1/bcV08rknXsJLmZd6T+4WVY7p6QvtUMcCDNnXOpvoGAam1gfhSKUiz/ebrXf7/TyIcraKNejHuxPUzCJE1YsgL8EQdFDiYUD/Exck
WixbdQJdBCTdGUs6SfB13acdf0O0RbyzP/17EhhnBKd+l2rbuytKyd55dcRQO1un8leqH2zkEBQEyc8KTX6sTAs/sowXJbfKdzXLUSvjOh4UwWVADdGMkzKGg9rRwj9s
+D/CswDlcYQUYwREKX7gB27xbMZU4tkzt6fHUTD8kdtb3RKMsn0Q8uBOfI6ygeEWzGDJhtB/CmyvsI9n7NPASU7eV5MgXf2yNcbhTUmuLW6Bs6+IEQgEwoYXZJbv2z/o
qXFILwQFkgyZQUlNTA4iAADYKR3ZCpSI6lfMxeZglNdWtdTGtFi7fdXI4ysGTQbwlowmTY1LI6fNEQNOG5OWBA2eM3GI5vTUDXfoHQ3zOYVW8DqghSiPwaRKdGR8cXXF
yneIZTGrjETCai0Eb9CvTQBz975+6X1o7KGMmdlE/CdyqE7yqOHu5jPKkB+3gibSamzkXevj944nkhg90D4Mf3f2OwAVzlNpeOxwZWwn7uPJBHy8YWkqicnO4y0O328f
DRh5nLhw3wmucf5JdxDOFVce6iVruW2IbV1asqVYlN9/bgtDra/v/UaiHGoj5xkNCqfuZJqvMP+30lBB5OpL667ul+9fHIGPQo8uY3s/YovSnbeXrZVWRNU8o0zwuMbq
WnYgEER8Py/ENAKbWLba0FSbcJUZJeqv6LPJki2nTpBDwrqUhabUenTFibjM3HzreYNV6wWtjRZ5kZqIsRQyKT4BVl1Xv9yoDsv1c2UxbLKIfhYtXkXnsLb5OoDuDxRk
XICWHaATkRqC4BGGl4RC0vp+2O9TFq4BHIxcQ5sWspHyV+AKw3kPzao8LMediGLigpWi/O/T5Mb5RxSVDDRNp1yAlh2gE5EaguARhpeEQtJl9u3LFKCBCfiaen9qwgmv
82w4EaX7DfQ9sOfGneP7im+5l8CVVw6hGiZ8++xC//CdH3SS3JuxvWpt+SAqTGfvSrrfd03XDCWd/BXsUn1OVXLnhAwdoSdJC+GqXXMfl11vJAgfInpX8tW4Us10/y9W
/MX2vC59ZpkFA4bIzLQJ1eNqxVUQzdoOVwtllxHyKiU1Lsxk8fz4Q7pi74Tek4zzrSJTC2RDWtYVySL77xPckoUntmXz4EU3XSrJ5Dz+yIBvJAgfInpX8tW4Us10/y9W
/MX2vC59ZpkFA4bIzLQJ1eNqxVUQzdoOVwtllxHyKiU5+rUAz5DYEkZqsKwJJLmC9kGUZSKUs6nfi1sL0+8BFZr53+9EXAZBZucO84UTSXnbmcKv6tpzRVL6JwwNAYld
JryprLDsfWvjd9IOaMsRqJ45nbXifb/WIl5fHciARJxxVYjtUSL5PlLfEumdQlXK3InWccylkFdntcwVXrlkXT0AbYIZYO+Rj1ZZKtKzzdZUk8xtnfi2WtRkwCOlWQlx
41OfDqqZ79JIP8CmwBPGVZWRX7QrcSxPTG9QYvG0hxq4lKWUzfP/7M+zAE0cgjyva0kRPbjgKubnRcCbYBSHodCo5MKlboVlRIWPCsagzAAdObEqRxwpqsA1yZ9muzKQ
2iCskkxh5Mf7twcxcGhF61nIUShb8jwxEeS60MQ+pXakGW8kmVJUfmjT0npw1+Qfn6cgC03jFgWESdxecw9ip1+FPW80SMBiGj44uW/9++2yp/TZqx2P6f009kKNPpQm
bna6qC8C/fvxHNNWE0FCjR7rifXKWbttW6MMd2wNJPKP3llsqThIFpcFSH8ptvNNUH34NyzEKFt4WpX4qbn7hW+UyHfSox8viI08BbZFKvcoXa6AGH7MO6j1ImrM/IuQ
2arsgEEFOFtfjxghFEdVdJ/lLkJ0Ce6g01MAlLSqqyLxNNwJtAnhm2SgiFiSBDMKgjj7G/zdjypkzb+ltE0gBKMNF7TgRNCQDq+0OXsV+LlVHNEwjuO3tUV6m7vRGUty
G8L4eQn8mBA7OFuMkWrn3qRLUf1ynVp08mAKAnZaxYDMWWaeLtj5ReD3Dvs4LeIn9wUfL2LuSf0mk6xmYeE4SA1oJrktyqqKVW3rBsHgPKnzMYLDj6qAgIdlADn9Rwwe
W0yo93ShBIPz2US1S59yGauTBxN2TLG8/zfCRK5pRrek6RVk9eYdi7dg1l2szPIJQk9PtonLoFvZKpagE806oHHeclefU8DzuzuHjDndQSoqkbXQDkp/b/XwKifqGfAo
eYNV6wWtjRZ5kZqIsRQyKbnwPsnesDtpXnoGBKCW+/v4a0wnwz5ZMrH4SRi3IN5oApbIN8soNgcrUzH82JLRIZCoLQuqG3EFLEy9K39sSt8jcWlwlzegqyPkqfw8iNj8
LvMaJyGpSnFvoHZarGvIIjNPWQq0Ht9vNYIslqwUwzpQcmpff1hRq78onTDzJ/hjn9Kn7iyzahRMsT92P1IAMQBcHKkn6ywLM54evSGOIeiGoVe6n4sSHW+kNZhXukIt
bagn9ruUgZYh4KU3+V8U9GYH16Z5u9aFjPj8bygWaGZCG/Au5I5ekz225DcS03qPSR5OqN/CJe2VBiUKecNkg/JX4ArDeQ/Nqjwsx52IYuISiL9BvoakLnXt56cgY2lo
iH4WLV5F57C2+TqA7g8UZEXescWCe4VAp5As700xPIjLWrTu6cGIHYSo91MVn3i0/lfsJ8cR3796ZYw9iXcYSuf/BAJ/b9Iw2y+msHg7oftykAwFS2jcCHCt+KEaN4ev
Iz11im55bgMwkfGoyBRbHc1x+EVTMLvbPWfvFy4RR5Ipd1j1V3Ecg1yivPjrXbF4jb3sPvv/07J5GZ55kjaO3hw0ZPPXdmMzYREjVsO4tYKEB/be7Bpd2LB5SsHNlmIA
vbQkvIXNdCrhh4Yrtehl6+gZQVFlMOd2PKh+nZx+ltF5g1XrBa2NFnmRmoixFDIpPgFWXVe/3KgOy/VzZTFssoh+Fi1eReewtvk6gO4PFGRF3rHFgnuFQKeQLO9NMTyI
yP5ABgHg5W2JzbUnC8zQ8ynQx/+zQaEHJofpPnJvB2V/H7dqWEaB7+MiXcsbldGkvbQkvIXNdCrhh4Yrtehl62VVF5xJQ4t3kik4XG+95ciktDxONjFZgSgg9ozlMz0r
TND0IKyT2BqVheFDnmm++vEdBxVhpHk9P9Exa0ty0ZpDhBt8GHG8CdESqtbGK36niTIMmLDUHSr3Pk7GCScgaBDSe+zZITTkp6NylBvSk7oluZCS6C3uGrvg0f4AvqQa
FSQzLxGPEwzbnkV3HPNJWLU35lRDf1wTlOW7gbot9YhcDKO+Yzg2b1XMgXIoHP+gOQ8MaWxc5jSuFZ7i5LfDmUARjvKC3x64hN+rnWoUU+qJYfPBPg4bnX3BWRMuUmhF
pZys7omTBktGWcZXa3mGLCfJwCteUJiUFB6IcCwJW/BEr6uV0U4PYNHzemdlapnJYhal3LeVfcGpbiny8l75eqNel09nGzm7BcrzgzfEDcQBsX4LnpYlP/OZ0DADTrPT
BSTta4dl+u+qolzKk1xBseXrwzmlFvGsW/pTt5C7zsO7b8Skrh8pA1jtygAqvltuoipuQFyhjF0iANUqOuas9ro5TRjQcT2XEqIRQJIzeFjn+SJUktM7+jUUOsyGwN+T
Z8AC3H3+ca2slGgSzF9AdEZYg9KB4KKMLjhfU3PcEXnaIKySTGHkx/u3BzFwaEXrztOg7Zp7iU71uDQjK0EjYW2XTpYP5W1IdrftZ5LPVFxiC53Z6skDl7GDt67YZKmB
B01TpEy2s/a7aShe8ZXFP3kTrMZx0KmObdQBolrUUBYpMv8+aZDlTgbcGYFsnfe88UHj/G5LaiY66pSBoISY4wqQu10KqWpGMUqy7ccFY/skzhRb08JkYbS1OseDcLS2
WFYwN/J/wB+C8MA9nso3Imc61MUaKFbvun8tXloBXCx0Z1GMqGPcgNFUBx+r/dz1G0810JlqrSPjLsRKwfYzlL3KLc5VkBJFBXFjiINZZGAhlkph19yYr4ee3iLuZA/U
FVnBqHwJd0AqlBHuxDrsWj6xf6SpVlB0eylLYi6eTu5vh8WMwOzDcoTNcqzDVf2gPO2oPqaDXSmfaH3V8/D7HCcyU1wjHfHm5RzRqEx90MXajmMEjKhUyEvrycEjvmp5
tq85M4qyW5YGD+EhLPHIVPPW/SPyvtDDde3gYkvzeDOIuCIX9+sEanXT937DYmS0eLLzAxtgA9j7F6cMHkg5PRuN/j0Z3bAWnzsQO3s1ddpZnFp8OXUi0NZ17JZS06uX
1TeX/IHbX4CIWkhBxHFUBidwzrL44cfL1REUVWFVHARfbORD5tWNW7cpEgh3qz490iiJlY9qNGNkWsJ6E+La2irCvJhoUuXMuPgYFodjJnp7JeJ2a2mf+/e9t/HOZi65
GECYPjxnbI3r0sFgWhZ3bbQ4cysAHmDUMWacTSDocPcApnXME6aFWfIMUCH2Zkuo7Ss7cx9wl4HuN0IcbV0BFCyJeWa1iDYXJJ5+vIfRK0vF8GmKz5YznKHq1g3JkbWG
eZ5dFf6SWFH1dEuM98MVtdxxdewatfUzEExvqDIMdVNiLOkCjlfJwWYHHaXb9+nQ6dDjYisAq6jzT2TAEi1muncPRcmqlqVZqeP/Z6PDtI+qNlVT2fS9B9c2Jx4TA0sL
opi8WKJjcV715cmhkVEXvGxtF70emwSynBRuVE2by6Q609lchZj671mN+6PusHiWYchSWjKJtQie9DcynpWGASMkjLEn4YZThZ1yQeFeyh4iH+CfTb1E8U89dykVlMJO
3HF17Bq19TMQTG+oMgx1U440iVZKG2u5J65XZRcCLoQAUVKhZ9poh6dvikyB2sm+yDRQWTGZGxOcRzXhG99DsBw5e7YDXT/ZS1aNB+hg5fSwl5RADBEZwwoXyW5sjrox
pPjGkBl2/lnNw9B8S8aoGHqCOheVsTmzQH0WK9rlux1cSw1A5W16S8hCxpwFCICm9PxdG1lU4rsCKdjJoZenqrdvFBE8Ge5IIikNReXdgZkXRbXIZUCJoLoYtMGXjt44
OOWySb19O2ZO+kszF/z5IFAGMNgewNK0Lh6RclDygBIe/qrOBgqpAeA+xeQRvOAxiWSQec8nTQGvhoRBg1/eJoSdj8vcZrWY8JoR+pvBBfImQWs2T0OyUM3WU/apzCuV
UAegqHMqXpWdFlO1xfrzNUfUTyJMEKt1bhKPfmtNw65bjRscSkJL9g+eyojp0ne01g3JHGUK1Npggc7Dxtxj4S4R/+gq3CPzh/3ZpKylosIaVPe+lI4rm3Qua/FCsUNT
RuLm/kxHwMS9lVf+XvQIqPzrjfKIa1BCQMJAhdx1Wht7XtQzGtpkxGxB+1LVIa5Iek6BSOMowEDzJ88geya9YEmFOVBiOk6GT2Lg2HMfGG+TwzvpkVoT1gSP6Uu1kMrc
pxxwXA70+4H+wwiH2lbZLsypnrJPilSSlrXBCDb4kVxY6sNCwBrJXVvO/mbk8K0xQ4aqkgPAxwQBYn1ufy17kocwO6aa7nPWVrl9hUU6EgiTArk4He0M7NsCy0tlUdhV
W1fWebjkkQoopBjcoG8PesGaJA3wCyLFfHmE51UJlAZ2qAROgCpR6KFe0uaAWTxlkQBtDhBpR6vs1hxSHAJjqSZmM438liNXlE0CjUowfopDICYq9+1p55aHzfiyzkrM
Yhal3LeVfcGpbiny8l75enqFR/j5xvApcZr2aGHBnggAeTf/oxOz0bLmcC2Hi/N76BggsyD1n/R8bhNoDkMRQAo2B0gPMGvIAoD0mw6oSDAJ3BDev2PW0QsebUtl3SM7
PugufUNA5DPHx5IdHR+CBW7jzqKSVOypZI4uc2W7spljcSuwwEfG8/jc26z3Cu1XmOXHj2AhRgh8ETYk9O7Oacc2Wv2ceRYpPSaFF/1TWMdTN0iCw2VQLcysmxK5h8mZ
ttMWzRiMyT/7EYt5z3csVoV4NeZA2PqN1UG8p8MBtqRZRJmXUVdLDrBBcEQYDlfIJskXu262fE7wQ8r4piCyjq8YlqUsSfDypUd19BCnHXnq2e0DH66LByVi3yf1QWtn
UDOtMMJmnONiNCZ3ouJTqmUQYga+2Ur3hlKIcG/nv8ecAIijwq0wfEGYRYFWLkunucyN40a35TXix5Un+gtJHVkks0BEUNayClRcXd/LksmyaWWxyR+zwqc48ix4oo0H
MbP/4aCfOb+oXtDl0j/dASuuCmXykb8aeMIMZ2RBZWTcMJ4lQtANeRBnzze6avyC6tntAx+uiwclYt8n9UFrZ4roQU7D2xn68KSVhAF+CxqmAMaBQSTUynyFmvmK5Lk6
Wl1vqVqyOnRBdLWUJmYiWmjYAGgKMruYoED8tHJH9eO2gwTd9baDJyHzY89omGucJPebLEV6XXzgoga/XZzf+f5mtFPyYHpBC/dc9q6Lgc2mAMaBQSTUynyFmvmK5Lk6
DZOOopf+w2zVQxC0n9NGNiNbRMcWa7ReHA0efWt+H90Qcsi0fci5nyNJmBkwtEpKSPvVIC8ChL9mR8Z+tUanQbbTFs0YjMk/+xGLec93LFai5/7dZy70tq4+XB5xtWcX
Gr6rM/CxwuXoNMGTf6nbbDuObyW2a8krZYjJ2TQYhwEBNK3bYYOzNi7+aJYcHHxC1gYMhpPK1T0ro1rQP3BBu7ZZf1POwe4zS7D7hs67n1SkruPTwH9SrGFunYhzkFY9
qQmSbwXUGZuBmaLevh11fVN/yp4qFCym9EBiKfry7f+S8ONvlQ/kGua9tzhvqgk8PhGk8UdbCQxoBv8rJYHjcdYGDIaTytU9K6Na0D9wQbtbh6F0O1vFZP8PMhi+rzgl
hB90RqAUo1HmxiBXPmut5DZujPngOazsf7pw/b/vT2EEPIQC8EJTbCvLgpP9brm26tntAx+uiwclYt8n9UFrZ86dNOO4n01Y66tbcbxuziV0VbtQ6iaPfXGE4c2/8J7o
pSnTo2rsBrD2j3jqfESKaHYkmgSi3odG7s1FWyP78dYxs//hoJ85v6he0OXSP90B9vJIX5qQ9giXGbl+k/8ml3bkZkpPbQQLO9ui2Cb+C54dg5sWs3VWEa5vGnpFF61c
nRU15HMgzq7NZtWpBo+xCQNtPNvbKUUEP7j7ztHFZwAxs//hoJ85v6he0OXSP90BPqXIWNwNLrW49+e9D5yloC3uLL5IqmSlJO9Z0L4GNSPMCcOZ5VKQgQA7JwxYZ8Bc
a9rvGLEkZj0sNo6ghwDUWWzQ69BxP+Bci9PfpzhJX0erw9qUoaEBk3aTec3v69bkYhal3LeVfcGpbiny8l75ejzdHvH1e3ZrfR7lsGQybiehex9PcS/OdjmLHLbPPx/F
8IHb8gzixYVP5O3QOFqivKN/c63v04/tCrDyYxXz4r94bRz2UwwXSOVT1DFahR6fvvXiYRaXx5mcM/DPkP+pFLE+jsuWak5GZUnpxjbwGHa8oUP6CDmMCAvansHFFG3/
zkAzW589VGPd0hT+FA/jT+l6p2n3JlRPC66OGCDhs3dW+SnhgRSJUv8zCc2KdIYRttMWzRiMyT/7EYt5z3csVjc+8oX9Q/b1Kc/SC6zUOdnL5qy3t1SYFvSHxJkEPvZn
HYObFrN1VhGubxp6RRetXAIqQw5leM87BVfc0NYX04j3GOXqeXJnmtMWmrJAzlB98DafdXZeXDCnTBSEct6Lp37G2FfOX50Ixz+O3ggHtd2HPHAcd27kBoDyUj9JHSlG
MDOZx9mZZIqrZjnWBHlMgRyipIApbGTwtrfHm2x/EXiw0xUr6QGQi8FNZZAJ1GrRrBIFZrIp7hsOyJva31ugR6eBKoCkTlOb1pOYpfyyTa7zgvQ8j/hGpFDEzGzO7puV
WowXd8AnUFE4RGQxALE9e4+EBz3qzTbZDR6VUSHl8SeGcQVx10o2VPg6yw31UMLz7h7zsdE7Cal45u9IR+yDhg+rnG858LQ1rvL+p32kC0C1MpkZah+hk3TzcfTShV0F
hBZBmUUFbRE2NMdt5sO9WTkqswDDWc8kTem6V8gS0qUwwLmzXEipMGloH3SYPXDkBhUAjRto1mGX1Ctp+dg+kOPC8sMIYgwV7l2+9J7JhTRGEu4qh8Z2iu8aUJKAQh1T
z/Y1QQRCBsdkiRxpsL6LyUtC7jeALL4hlAARpHYXZNDlcsc6waytpevht/IYEC2tHxwZkg1ukIzeORVORpMUv3SJ535p2nowwxjFrN9vw9rDszeJO2Q2bgmgu/trCr6K
HklUksmBvtBkHrWEoAbZ/HFtywFR0S1U73p9jpq0GKIChm64ayuzFVbzO6Fw+SfSv7TCsHApdA6oCvaVwNx/kIxR5EmNdNsBep25R3GmxBkiST0V33ozjr/jrvjTrMFW
0N5M+1NduKB2zczhPEJjeiB6K1ZU0gAvdoiGGbVCw6p3EC0SmkIMQOXtsZBt1G/D9qnntsGroJYNHfV5yRpIh1G8ALJjXz2FQZ93P8eMAo5kIJ1NRFn/57Sox3JK6jFN
vgj+Pjizq231DvfwJzYJ5u/QBWqZ+McBnk2LgVX0H3i6ODqUQ0YIvPISHPnPfW9JrjnG9x2SroW54sOuUlxm0y36RSEeHNUdS7mVvlbeHovh1J/copGZoGTu/mW2vP0Z
lPTqS3H4GLPJzAPg6u0iKu2lTm3O6NOKJwOEJ7NZjNM7s0JQxH1wvYsDgZ+pR8m/Z35L7G+348aPPKHhOg2532HjViqE2rAXPRufnkvhk6/NFdpPQWk76kYNsyKk068F
VrCEYmbXhpEmlgx8prFCF8fQE725kM+r/mXtMkCwc3b5uAhKbX4zuztlIyH4ux60s9gPTB/G9nu+dRO8ONuT+CCd5ZzXTepuJAdfmLHvrCkR+YWp9P37wXyrZcqIMPcP
PURo/7G61bLbg1WaaqR2XxVrc9Qx6uLLj4CQtt4QJcyEwHuk4g+6erNffUAtMzT/GjLGpQCeoSf8pH2DEGFmEzET7vLblXIlRioXOf5YyF/td+IS6g0W6kSDE0UAGx8D
VGsBukEADrlDTFlWJkDklV5AhPzMSIlK7ul799XlnblLbAUhSmko7c75bIUl3scAOaccg9fUV2jsNHswv7dbx1DqhRfsE/gHcsKvenjy8R48v4RMj7jX3BbodRteEr5d
DmfN1LdmGrfZGz/7esO48FgHDlZY0f7z3Os0UYK4WrgWVNVqIayEp3+00ybxK9h+chP4CqY2MgV6bRT60HUqBw5Oj+pvFRlXeJC3RrkF7lFML/qarIhzXb0b2R69CnNq
gkQrAa4f4DgawGJH5wdgPf8nArhwIWyPxriQSY/RUn18FlJsCYQZRcX1ePvMnb5F7ONpTej3iTc1GKHVp96MCLaOGZL5L3WZT2WL68DBKzaulT7zW5acpwmy2Qfo0waY
VchLOMD+ssvRfBVWZrRtFH6A2j0uDjaF4XZviQq4MZNRMkyWM9YkJ4Xn9YFMLg/qmHodDwJEgXidUKD2RaHh5SqsJ/XndQd7AemEW6vp16S2gwTd9baDJyHzY89omGuc
C4OnWxQBtozlOkhmGnS/OjFWkAX5yGaFRpoKI+dYdOA8AHb+Q2VZHXZxQwFOY9TW/uv447n8GbnsAIEr6i2Vew5XiVbtLiH5hprd2evLA4mitx5ViJsntCTUl/oL3Xn/
pW1P1XtPSGh3utJ44JTAx6yC5Xw4K5gttztiuzRCVFf/4coixRt6AjtZuh6LgP3+OhW9PCdDOf5ztS7bHKpeF6yC5Xw4K5gttztiuzRCVFdGLUuPWFDBNpZOKyxIv0jr
9xjl6nlyZ5rTFpqyQM5QfQTzCntqxwuOo0fVpwfjzKJRyXoGwdK1xExYDAnNZjjGC4OnWxQBtozlOkhmGnS/OkHj94M7aiQ5Wkwne6pR3IF2E1m4SnaUDZVtCzfPF8ey
+r2QJHaIbmNea/usnBZAjTsKy1ECJvI1c5mv9NxgZA3zus6mTvWkl3iV0s4CxQbOdFW7UOomj31xhOHNv/Ce6PqNz9peeAiz/2vQAddXx7UuMwysW1ZHsZUrXXlkPyIk
yM0Gj32OqI/9O3NT37wtTrBDUcQ+A9tuwnzHtzSLajz4eMNJryAkNGHNwbYxX1FcC/8cLDKgpLE+MAs3xZb8OIZ2xGaArqjbC8yQth7mP0M1ZOK3xuPlE+3K66TSI8/1
vHcL3e9V8Y9sSMU7B/trCAuDp1sUAbaM5TpIZhp0vzoWS5vIP0RT2SQXsmc2eu5SPAB2/kNlWR12cUMBTmPU1mR3yZ1AJ+aGbrAc11Jgy1eCll02/Tc/p2/oT80T1l69
khrXU9l2MCj4RYtQcdRVToQs+sX6YZ8VkKhwI5v97vYDOoaClO7v6hXtk4CT9s1dLhttSCm0HBI3cLOHI8irTh6BDq3KJo+JIUvrYUXN+GY8AHb+Q2VZHXZxQwFOY9TW
6XAoQqV9Fkyayq3Fmja0SsjNBo99jqiP/TtzU9+8LU6ZzjWJhZqjldOVYg8Be6j9ZRBiBr7ZSveGUohwb+e/xwef7LcdBtDRfjn8yCEqDtRH7aBI5f7m+NdczS0bjbxg
toME3fW2gych82PPaJhrnAuDp1sUAbaM5TpIZhp0vzp6IR5QuNkKmIZHydxxZlPls/Hm+Uf+4c3nUWQCiGg9e3/eofOt3AaedsnG61aCoz2EH3RGoBSjUebGIFc+a63k
SayHp7NQyBS8ARAhjcW7PYuV1K0R4eJgbSq7szcw6NpmxMkqYu+iqidhA7+ZldU+ejvboF8NeDfRmuK/dlbYCnm0MeIbCzN2fFsGXJNPjVXos+28aO2hajUgEcccp0k1
/sk7XprCPQsYniUmr/ycO1q1qYT5dqFuIMttyoIc06Aw2A6OEX/MFUVLSiPqrUI6f194HFyBTyRe8DdUcvoQ/dfcWe51lmPDHFHqVGRjYuACvCQCjEy+snual+IrPK0V
XI+5KwDAmf4Eyf5Cu9ZCFaOYtUVokc/l5V76477ajfa95/YQ/aY6rwuywcRqxvLnHNlPTdI8po5DL5xlvbNJNCXUJ2ydMqNXcK0tWH8wLO0kBstI1/ZbCv4r5C8a3Qrp
1P5rE79buksBPWaXJsufYttqrEFdc8am8X5ZZLH9ns99iUqju8aXlEUTtTTCYVXkOFiCo+j0w20J/j8yMIzUHroZC84Wm+ngSwFEbjg+3fTXc0QHgDZfmraI8yZQkTQf
AQnpQNSRgvXoRTy/rgqHmRPyI0FsO2mx+UNIQGk+FBBkkCIzxr5h1s75PXVrngH47FSJ7I1X4xrUEhJWv/Gw7H9uC0Otr+/9RqIcaiPnGQ2W1ydMHKqIXQaAiKeBNXkL
6veUGDef9ncH6a8C8g40LzG90FLaLubniVNhhV119EHUbOGfFXK5qGOT/immwDyRjhLPVzWGO2XF+CiTlZMYNVPCNzLgsVbBqoZK97V3YHcTMoSXybtUlLhYOQD5U857
2z2I48upCBC49eX9kgICzG/vef3kLjVTFhbmGIeIoj+NfL0qkSKE5WdS8jQlrhBezInXbV5Ue5TWkZpKiZKzpBpytfCogXr/X4GNlYMU587IZEjd4Q77rDtguwC9Bn/2
TiA3zvPWxafZwfHn8sVy5Zbvj99dFxZ0/pUqsjsVweWzD6MBYFAj+s8QxuvSUefjttMWzRiMyT/7EYt5z3csVjiloqWhjGXFjBTtmWcYNENx5yHXJPcd8tW0+DfJVt5i
A8qS2fXqx1s7elsdVGgPtTkpkO491FLuhBpqHxc/eTSXlDGS0xF56oz9/LlT76vgmdADXrSTYTGhI86chEoJGvaVES7qvvnPS/aWjQR9sHy20xbNGIzJP/sRi3nPdyxW
OKWipaGMZcWMFO2ZZxg0Q0OABU5jsZOq/oDygAh6JVGREIcJOi9AFtW61bxklZAxgQUJeTScOhywIA+smI3fMsWWPJWkLcjGjFe+Tk6rRYNIV8Yoss62IQEgUMTe7YKR
IHgHIbmxj4omSSy8PEkS+kOLFdEyhXqtPCPEcDCye1nG/e/WcdkE/y5Rh2NGJE1rPV9qh+LrL8FGC3cJw06rtXohFhg9IDBxUwOr/UKSYik+IfEzD0Zs/trnX8Rih8sD
uqZDxE9nmB67A2N4jaGr+ZLbcGIUrmy7wdU21T3BCNWmA+lofXo91C32YBoUQid16FGcMo3f62/H46i3zj1O0+sHKb8te/SyfQKlGDCevyxhyplVgxmf8NCX/auKfY5Q
OUmkFlmfNx870GGGL73aj9fcdNohP2x7PcPQWy+46FxHmAGPDvVT9y1EShV0F1Gn5MtAVC1WT4x85lSto9b5z8+uNYL6LUdxSt63zwLesrOKM/+hTUnLc0UQEyS2JRRu
UpzSO8GHggIxYU/n1grL/3PGzM91e/fbTLsrQg3nPQqaCFbZgurALH6uC4/JjhIcrf8l3CZzxsjmpbuEp53fQ5YiOQhuXG+GNDkWIWWfPVGpNz3BZyRTDSSx+/B1280v
z641gvotR3FK3rfPAt6ys/QseeKR2ACrTEAPwZ8IL1FD0boStO358d9NVRGDt5hM+1VE9GylsYfcBN6m7Qo6yMOF7/qDqwuwnYhI/F+nwspCxNcCJi4mih08pMktR2Ge
Mk1n3AWs+o2OWcINn/K5G1R9FtHjXD5yj+a1AJZ75rfDKySKb0zi2YNak0QlSZ0PDegG6UNZRAmT5/S9rzqUqmLnzLrUWgS+9oGs/106mixCJqI7poNN9SOJFYmy3LIL
rYeYKnMWHHHlJnkiDoB18RhJDFhTHBKcNvldRHCUtAv/DJ/rghzG9xFfyUQC47mT9iyM2ITYpjW/Rh3CxIGno4hYg58aJciIxinLlF0VzHBL5KfAoAY7gNDiOPr7We6a
ttMWzRiMyT/7EYt5z3csVvUqZF046OjdyiJHcAwKbNDoOny9hD95m0JB4xDOhPxrA8qS2fXqx1s7elsdVGgPtVkOR7M/oSuj6MdNXmBUTxPIZEjd4Q77rDtguwC9Bn/2
PEYX20+68LII/NA/VeN0OOr4E8ryaaSf8yql/rjrJiPWZofuWyfxD/uS4/GrEKix6tntAx+uiwclYt8n9UFrZyTaICFQixu2lNQp5yoqv5QM9LO5j4qUNZSCgw7c8Udt
DlRN8O18zQ0vsbsoDL3GntU6GhtvodYSURtsRMet/JKY5F2XoQhgyzgOkhUlqxqzOH9l/HqczxQZlpeyMv6CkB9ySK8elbJZonwJmJNrdbZTf8qeKhQspvRAYin68u3/
fU8Zg2x42Savm5628IxG6mygsT6uRkvKnGBF52nc/pVXAJLMMwW1xPXQGIwG22B7wHn69TlAn4yTCUN5AkakTLbTFs0YjMk/+xGLec93LFbaE1nb0fR5maCBCgTY0LpO
C81h6W30C8rVTJEVeAPQaMPCl7mRMAUviJbY1LXDaYAh5lbJabHJAbgpddL2pQLbyGRI3eEO+6w7YLsAvQZ/9pOkraUhKO6agUQMOMVkPnvzfHSG/ttndaRkbjZYts2b
kgHu1YmurpIMGsHMh3fYbscNzglwnwzWyO31bJjKyIu6pkPET2eYHrsDY3iNoav5IipuFwAIKX7CUSYqCb/fcCuw7+pLycEuYSl8+neZfTJ7/o5AAS+3IW0QDUqXfber
GLY+YSQvel4ENa6XuaP4IIxddXAEwnGrORwH5/YXUy1PyjoKYrqSgdDSmzt0G6fbG6qyqwXk5cKhMIiKig7xidH6UcOuDUVUB8ThW9EsSIao3thgYWss5afXiO1MBKxh
APx2SV2gDnznnFUO2ymoyRUp9kfxAqJdd5GgM2t1SxmfKqhwyjTQUdhS4gACW49WFUTwMIFsgiPyLuUBFZbhBcf8WGkbRCoA9BZ38dXyWwVf2MZ5gakHdTRH4SE1zxE/
SlP1Q2MnUEckpvskY9PJ44MQPsuBJNsPyFGc/rKqjMpC/Oor2y27Us93O+sv4Q4I6X1SU2X/u1RJEi8QgY0J7chkSN3hDvusO2C7AL0Gf/anTBDfPC+OYLsfNqQKQxhU
mPOoRzSdnCTm1/CVCzipZQFK6I8EuC0XejwNfaAHIdTSZe3tscisq0EtywJCMT1flGdwlSDLqwl8gPwUuzxbVFHtr4fQQR+CerpRBuHZYyUwBm9i2Bpys10uAEPP7NPr
O+TOk2uFSHn25syWL1WIsyBmHmKHYdsuVtYkRF/aPFL7VUT0bKWxh9wE3qbtCjrIJbW/atUMHz5A1jZGIwciFfmjmgQRFzZU1HJl8NB4xC0BiD6T9DRWR6pr1fwQ+r+b
lw29YUO8rwK57OmSVuCGUiVpKWMe5mOL1IGox/M6AgOd0kN7Ls5HBQ0iMqqaPE0HZIIuvHtXjX9pgEWoJUhymWUQZu/Bo+bRqT9CLcAXzUfL6l0W/CApcwGsXW9k/jLX
rjhT4/pgQ7qhnrDTqnGgxJluZscmfuve5TqVX+l9+PdUk7SkInTJkVQsgZsUYF+cLmRkyKX/JG0he5NptwqozWz1BpuhEgI3y6gL6nXp1M2SrRzMGICL4LN0PkfuqgKf
q3Sa47bTrGgA4mOjOT3Rr/2KaoENth90VL9Zy2JDreSRcta0D9Kj/VmGBm+qa4X6bJ0g86zc5qOAs+5J4chyGw/zxvkLSiMyv/AgsYE6K3bVbyQ7TFbPF2CK5125AeXY
vZEgSExh/6O74WAqQWkc5yjElnmfScrhY7ed+egkMnFpXfJ8ibt9B7mJXn4ytASvw8nrsZ2kFDdy/iUmHDm220+KDGTE/fn8FvmnlD/ZBNNCfyK9stBj9B3DzKQsg+Hi
nM/M7Geqx8qUWQRtRcJ7tZRncJUgy6sJfID8FLs8W1Qe34koFCJZFqp4GHr4tjKZyGk7KRFkk4Q5fb/4Q0aIkYG0lVeHnpPIrm2FiuED2XMRbT0N8mJHwvDXBuuNuzum
QNTocEL0Jt8xajr+zIYT/8rlh6PO5G1rd1rOQe1bOhD/zDiar8oZbH/yI6IHJJfQYJxBC6mUHyV659AQlrwSYMBZlG0BNQib7IHW/yojxUVmQTv1/L8bmpR+v1xo1TBN
JDbsOKebu1NdSu5LV6pANtogrJJMYeTH+7cHMXBoReuyRbMSfoHhbEFzTNJLe1A+xjynOuzN2R8ibxRighP9uSdRAj7BTWGmx+/yxyVjb+QT+d1XOXsRNUeYL05GyPrz
3mAwoYGvQzMEA5GAEnetRtiqesazBJOv4pYyYFt1LHz+13+HYSHNjBdnS40dss+5ZYZ0JR94hGOiwI5Ug9uAICw+32CVi+O6DYx6uGbxQA8I1xtDB6oCi63XMTENVpnp
CgOceyaOb6xEYFGqYrwT64f0L1xgMgEUdTpzipGXIXAFzfqEmtpa9jMjGuzfuJcCyGRI3eEO+6w7YLsAvQZ/9g186hXSKqh+pbz7VnwfKs8Z1v/vl70R8DrpMeGOtStb
JtYNHQBOb6oqNemXZrG/IMYu1UYtFIXk2yz7AAdhwWW6pkPET2eYHrsDY3iNoav5dxob/wuG6etPVjyyTgLH/Knho6G4QOMWMo9ar3+1+YA+1Uyq/31D3g8ZyKA0/wJa
hQ99vO7NS/rba7iBYKjh2TRF++T2Wm8p08xaHmzk1O6x3Y0EIwr7vToCQrFtxAivgWOA4aItEG53O/F7OqJ/uaS9qFa0RHiL/WuglJga/bYlu0RrqO8D4F7gL8hfEu67
XAYZwlvyyYkg3Q/X+FIntX57I00W6mWwtSpKpNmmZM8vijAYRsf5XvZjAkVhmA+Nz641gvotR3FK3rfPAt6ysyVB6fqn1VcSZmT0DOxQ+B67mAdG8SYeb2pjuOuYj6zr
jVKTmdYaxIfw9J12z3kxW2HKmVWDGZ/w0Jf9q4p9jlBkQ3JyVgMG+XJtQV3nMjYKw8xt330xBrmkfwoYy9Ihr/owlZ3Q4fMznQXN8GzGPDKaPloHFGwCM2EYH1PrloAM
SfAyPugOlWx46j7aFk2+9yuVhxmrgXPoS14IVfgVcMq1fAe7NECHzTsBXPzJPsiwh2/IHQ3eZV8CPF07p9087ya9wCSVG6/XmXJ64KQtBqtWEMRl/JmbGds8kEst+lap
Yetd0zYBHmCGtMl3sGqR0UkUTqUtY93JsK0FUi9FS3gyM+VXGPxsoswnq9p/+nYZzY4kzgetb3aGsn6l7P3hqkL86ivbLbtSz3c76y/hDgjJPc8djYeIqlsYd/aaIGLf
AkRENF67A0+U8aLZih9ajs5bRduYDDOcLr3QBTazFZCGcvhYvgnPXOocA3HALoWsp7BLRceb5roF7+lz2Yu/n4oy9BdaJgXlRuhDhj2LHGGCcir9LqgdX/0kyoEJOe88
jjr//Bs2ih+Um/XNhp88bW5F+kIWWu9/1dFQLvuwHL1o9baxXmaVnBcIf2WciKpR13MJlhY1TM+RrMO/+ix00l0wzJyYLf1g44/USMgFSaO5mmZKWW1U7YeLJJCCa9FH
BcsjjdjsyfmBAOCN6o7Qa7VcMtZe7r1NZFPK6gCe1ETg1EUWBhAi1SV8J1C+emznuqZDxE9nmB67A2N4jaGr+auZbl3C6arPqloTwKtG+x99KjaW0K52hFGM8TO9+Ed0
W7M+RJamIpFNXP8ok6QRlurZ7QMfrosHJWLfJ/VBa2elS0aVqfSsILg3azZRu2+I5uLeb2BA0Q/dLXBPk+N3mE3I+L93kaW9TyNKii1rU8hhYwgvsoOyoX653BeDsZOI
KBE4kIGdGxnXggNWr6Vy9rCukYDkjpthmwJHlwo4RCEVKfZH8QKiXXeRoDNrdUsZBgdVv9Rb/INWOOaOFKA2ZSxY9Hvga7IPzuvx7x7wdciXQ/e0d0fQYjkqHlu3qijW
cgnpZPm9XStiSpITTNpoOfFasIj6Ev7IHC5sCie6NUbdImymrv96Z5+0+uWIZTSo+lf0OxvjX5eanClUom2DMyAfqr7TKHYUB790V/PMU5YIq90FtRVReggkQn0vvazK
DfpttSCdjkZKSdACLPpN2HCHx12Ppg0lQA6G6QYBxCTeqCMuGCnTbfFJZPCVb3T/hRu9XRbT+Bf6Iy5LSgaKe34UeOlgmD8qRY3hLiZyksu6pkPET2eYHrsDY3iNoav5
4TVRZiS/7PGFw4EbPiRGXgp6VuaZjJ8OJ5DVz6ahaODpDKPEys1zPSzCsh9HzHPuhQ99vO7NS/rba7iBYKjh2UYUHbdWljQgwfTgcoAqoiwu0UJ1cy1thkwCRPqmYQV6
6BBsBSdfoadzT9YcO7KudO70d3UQEzxqGeXllC3Tfbq6pkPET2eYHrsDY3iNoav5plvH4hICAslhjLiT9Slrc5LgElgnPjvpNaTFzGmkl0o4oIWuO7QQpp5/CEEjneE2
0l7YefpmLImuIM6RskR0RSGrcA4yq7kzaWyR6QW1tYw/6l0MxJux9maJjAQL4sAxJWsmNlPZ6yDqesE2jwQcHYUPfbzuzUv622u4gWCo4dnoO/ZUo0T9BiED+ABG8qi3
wbygsjHs1Q6RgxtPtic3DmAuyN6J/RNUFSLBgGVmYjLwwO4kSFQo3cfX4i4M3dUTnNc5FjAOqqvKRWwITNIUsTrQ5oSr3SVGoNzcEDYOcdt4c5QzMl5oAljqUh603nnm
AuihlyI7GPxU6xRHz+T5TGl+OmWTgOcZ8TqPTXqtiu6HcJZX/QYds7vj5AaUb1tg9sLHg45cypYsX5TJ3KBZnQrFsbXO7CL8sWgBgJU1GbNzrb3yMrPANK9l+MNtewWC
OUKDSbctgVvOOm9G9bC1RG30ZrZbhkRqjCCrIHtHyBsE4mDYtJV03BpiNZxnTJpvn7H4Dome2k/gOmpRxLYw9GhthetNB+wBxMMG/+fKlUklaSljHuZji9SBqMfzOgID
gRX616DtZXCN/LPoATZMzwi2VmeD4x1a0Q41clsteSW0XHzZRS6PIAYpAq/2nFbhOb8sBapoxBfE0rrIGsVUj+rZ7QMfrosHJWLfJ/VBa2enK+7OrC9JfFlWNkYd5BQG
lbJlzhwZ/cmRUG1A3hemOfnMuP6gabvxpMBniTyRIZ4n1hBBlNR4BPlo0ciCIzlEEO2mPq1K3jpo3AYaAKPz2MY0JOgRJW1+j1emdH97noX2PqLEjwI6uj955Cv6Hcqu
d1Jva3yRyzFSjiicqTsKl4rWm4uhpGmiq90y6IZhOaXK2KVyvGo0N22mbVGWyj6M6tntAx+uiwclYt8n9UFrZyYAp3d6zByuHJUWCxezbO2VsmXOHBn9yZFQbUDeF6Y5
imPqFe1F/fdE0ComRFqeexMX1IKCfTOkAgg+HM8HBJgKo8IQEbs0mVkTPALSXgvKYlaNYX6bsz32e1MqZzDaup2LF1W033VC4N4FmjVOzy9YSKZQcgU37hRJ4NAGTe4J
rCuysmWPcDG7Dv5jBMVDVh8zEpO5O1icxlwtrl9SX2drfYX2daRSDk5+40eQ82EboPSao3XEvqB6AvPISuA90d2SI3Uwvrs2ricWbnHP/bOhzhXsoLEpPJD743j6y3JT
ArjS7N81BCcY8OjdJeAFamZNbP8jHEjamxUD92m8ZCbVqTBflfxXd1etNMte0dRGO5NKvhzEnJcDGTYci1pM9ihFQt9LAcHNdCZJqB2AhiAzW7dGR0/PkY/V/wyznZlV
fdIs6u6P05Rg3QNbOdmQwcVc76kbgsgdjIXwq1oyVELXAWs30N0eppPnvX3gwtfyv2guyQcoK/LsGK9TV1e6HViZShdQEbmrPDrou19eh6G1ME0NonlnKEx/uQin2axo
n3AlyQNF3iH9bLhKdTVveRhJDFhTHBKcNvldRHCUtAvUJUCpdmBOcLaGW7juy+5NVriOkyV3xeex1embQgq5cnohRc++G4gsY/sbcV4dQHjNpKGsd5QNtYtZ1dBiXWdx
HYObFrN1VhGubxp6RRetXOqBYu2nzKEo7CWT+9rMki9IDlpC3sj1l0rjMZerH5nAYB0bf9su9XQQZNVd77zRMOPjE/OdWBTyw2La/efg9aWwzvXk+lWMJAnLOpRauDOG
VEUVdMD/Vf6Z7Lxalkf90ZRncJUgy6sJfID8FLs8W1QzxbBvapyVDA0pESgvDsPUVCAuxUVvchiJN0F/46nAZrX1vgUq9knJICermo5DNU4louWIisQqB3V6AdtBoH1K
PrYDZQs6KfAuf89QV/umHcbcpxBMUudf1NlaZ9AEXHoGLtoHB17DS4HxackxeDsE5aTKmLttbDAcJzy4qE53Z7qmQ8RPZ5geuwNjeI2hq/leHZr1/H4b3/4QWqkW/LgO
Y+hbuMDLq9BSS+8xd3jRo2VudK20oWDkXiRO24+dbv2N4yy9LM5PhsWMeLUHMubbfNPkPLBbkgDLPqaqdU/8XubBQng2z3q4BRyb/lBiy67mIsbdrGNJL8M0I2PA7PTl
gMbxwq84b0yzt8MkWVTTN9JqZhMMGDsGEenItHZi7fShnwQptGJ0ffnTvbDjsef9hIDXNYuRbfl94vcCiVbr4OCYpDUfRQ1NjSooOjAq7iz3l261tMkyytAWSlvtEZUi
fXgScdx/u3cPnvxXpF7t0gHhcXNTnvWNFNZqJ5PPALml8W2k7VvjQGdj9RgIwKkyuHI4IdqbgoWKs8IW6R7N03GZnR910QRR1zBZ2R9iMk+iAAsuKrJ5CQk5xJ35wBcU
0fpRw64NRVQHxOFb0SxIhouNqQvQhAw6jI8IC5ao+MOkhWQZZN9ZRsDzNidwcaOyr60/fgmNRJkdqp/U1+qoQQTaSNwcJDS0zxqAAHVskJNIeg0lprBr1rDtef2shTsj
idI104Vxhj5wD886RL/XrnzVQEToEmYs9WztJSzqZtHCxHzBd1FeZ4LlzXbbPpSU8UEPPsCqAMlnzaxIxboSFE/rf91JafTmVIo6y1lJ6TLSECwXDqwXrKSs89d+90M0
aV3yfIm7fQe5iV5+MrQEr2nsviqpMtEaTahAYNG4eOCgBw6nZpLo5jLfP3pdhBbCyKP0IuqoDJqrv2dkIPx1tPQiIIFXR6T385ccy8whQPbPrjWC+i1HcUret88C3rKz
2fDqxDNUAYOiPgteOHRKuSPVN8zUSCDzJb2Di+Dxzb3vEOnAvK+8Sfy+DuLH2MjairC5OU0Enxuf5ROkS3YcS/lvcAfpzmbkxrZO96HuacXBkUGEIOpFN7UwmzBGJQAp
ttMWzRiMyT/7EYt5z3csViwdocXLoIZb6euMipqtrC8hL7qmXBTUWXfEIogPpza5dSTIF+tlRnnwVyIWy16KIyZ/VJB2mwpRzV9WBYjTwqKFD3287s1L+ttruIFgqOHZ
2a0SNMON4R7OMRcBS4/dtdG0bxwI1G9FwdYV78j7L99gLsjeif0TVBUiwYBlZmIy/+oNDz/XIc+wJz/oW4U1oSW7RGuo7wPgXuAvyF8S7rsCiq4pZzKhgle8y3FJDqf8
Mgr5T8mu872m8FGOvhnkup1UMEpXkzM6RsOnbd3Nvb8laSljHuZji9SBqMfzOgIDoJgsNzvtED/9lqYjXEp+yqUXF+YK7XqlTBxZ6X81HDA8J55jEqV+4X56HOmjBO4d
P7OMCLHcLlHNqe3+T7Hg7+rZ7QMfrosHJWLfJ/VBa2fEHwElk7rn8prH7PTgeXxtXOEtuklgefqGTIXpoob9l8CJ1uPFT+/itpojVW0b4F/tNVNGGDv67KQSxVer0gv/
Mk/8S3sQNtKYSfRuBc4tBEnIZ8afJdQCsK4G4hG16VR1TNFkBRVu4KZrQel5xf2Qm4WzcKJCjX0ViEbR2pZlfbqmQ8RPZ5geuwNjeI2hq/mPqr8tf+B6u1RGltkHk3ry
CnviaRMvF6pBgmshTO2L1k2wVM7XcxVsUh0xuTTKCLL+jMnk4Sq0XSUzpP6LaE4AYcqZVYMZn/DQl/2rin2OUOBFjKQoILx/uYlAigl1hxnQ8M/6eyvFUEV2If4tU1AD
cVDK3PQnMda51D4MjJaGD7bTFs0YjMk/+xGLec93LFYPagn87F5P1dGh06gezvEeIn2kf5wJZqgUTsQKylYb57IBpHS/F4hVPx31WnQgkySZhwxypPQVKo2PI+K6/ZNK
0hC1oQt9cfCwUpPBqzdMlWZj68g6CuQosPSHLZbV6QMBoivC3U771kd2mPyBn0yPsviGnMhYtNNyhCKfWLN/ZC4xbNQB/kiwvgdtf73WBgnaV7Y7MuzBykF8JUWjpy3l
DGk/gvi1uaJKAk5v/eVngy0TzgcT3KRB4KLYF84Ml304YVKPQ3CFpV3KboQB9QC82nw6SxQVc7X8dDev7fn7ysLqnZTkTuQ72cd+riRHXPUSBsNepJXfIJj3swvh2o0K
scFmlzft46fzRBaNcbxfIJ5dBmlngHTGiWe3UiN4oHnTX2+4ttm+opB/u9DSWyeCM3UIX9c9+NTJ6SRJEgNjAC1+bfIFFX1bLUpJoGaJOGgr0KbpmTjT5lXcFY/3ZsD3
aV3yfIm7fQe5iV5+MrQEr+nYZkLxcnc7CXpPSEBBUVIT9vqZ+d/V4XU23j0laV9myKP0IuqoDJqrv2dkIPx1tE3n8kNTD+9MrNo5EDR/WVCUZ3CVIMurCXyA/BS7PFtU
GNKMpoB+GClb2XpvloEQEBP/DTdTA0dK5Z44vomzzYmEzGojTTk954AqF3QIMqhw2B3oUr9Lb2CHUltiguPMVI46//wbNooflJv1zYafPG0BfCw/ABr+f8aEAPqilySG
Dp1oPLAk2Q5jiirSeUgmnEPzJ7AhYNPDRfr2IUy4ZYFjMdPHHkxccznF+QFwVYdEQhBFiTcDLyAO6zValIVofdNcxu/yNTPEUKgFIXNUKptlhnQlH3iEY6LAjlSD24Ag
DarhoRJJCplZaSqV7RjWrQCOv4xM23QiJ82JDKKU81j9VVpDITja6tFKFOccMpQyh/QvXGAyARR1OnOKkZchcDHNLjEYRea1S5Lk9VnQf2Elu0RrqO8D4F7gL8hfEu67
y5SQjHm7NHkUTpy3QnOzu0ELOIkSNInIyaySwT2Kc4yjkxOA75foCpPpYOEBKBXjnSc8vVvlu4Cu4qoeaJ3p50IiDbXzcuAE1PuAB4AsYJIcS0bg8pQXvrmjZsVNT/vm
ttMWzRiMyT/7EYt5z3csVncd8fVwnc2YpjtK3mk5B7sZaHf2KNjcOrkslvWK+uHSCFy/hyJN71QJ25xmGkS+DtH1qrx6CtmLBVY6F7oSTs3x3XkZ/m+XDHl+Wvo2YzH8
qSiZXw1eHl5SyGbzC7H4so9shlOTCjqCvLH7e3Mfq/A9ZZkhyHerCGd+RpOWSxxzniFSVgNIQzheMm7Jp1ICvzQUkD+lyoh6yjyjG9TBVeLZ+wFj3szSBuOZ2+yTy3jL
ejLsCPAK7bJCoFkk8Sbzk5vmvGDcli8OzJtHYmSFd7bkzWGxlymbS/sSpWZnZV6aeokkYbop6NBftPCRfizF2SdHBY5nxbsCRQiLJ7Un6NTiK/7L3+SnZjbB9OTf0Z/2
uqZDxE9nmB67A2N4jaGr+YIakLQXPZ5lBCVawzPYYjeZpHvUoQVulq9+UU3WiONEeR7v/kLvltPcpwkYNgUGKx0Pg7GKe5l2a5Bl5NqCgjGUZ3CVIMurCXyA/BS7PFtU
rd9HF1Djp4QRLjH6121pt4NGQUE+bFnIk9VeqQTgJdMODFQ1nif2kQmXAarEM+9q2B3oUr9Lb2CHUltiguPMVI46//wbNooflJv1zYafPG1rPE73A9p6+c3jGwhcoHzj
eJtFD2/WM9nUAYLwCFcAT81xjDI9E0dYbbWztNLkX3UtV8nYo8apfyVUzRUxld5qVKPtx2VQaP9Ptln6+6MVgs+uNYL6LUdxSt63zwLesrPHu5vPVQq0VIxatmVgeyGn
lbJlzhwZ/cmRUG1A3hemOWATxHTdxb+S3ZHbPIRQLv1hyplVgxmf8NCX/auKfY5Qg6xgJQBBR2RbjvFd1A1HhDHqtst/W07p1KSU91jnTqBz+TITcMWVFvZzldIRXlZA
T7tl/YZrngvQygMs7leT0PUXrLW7PKSCasJzesxQ1NZgDaJhTEQMPkPPv8XzYPXS6m9BXH50ZtqcslU7/gfRrOcXp1TGLaWdIPx8IvGqvEEFSFQqf964k5xa4ysEokiB
koDBCfU289rRffGz2JBnz9+FZgozy98BwRZgddFYergcmxq3N/gPdV+unbwr5XWEmYSnwiqLJhcpbU8V+iStqdxnY2pUv4gZI44pmCGR4ogd3sI/ybKcldQK8ADb9SRz
1pNGdeu3/wOtFOcNqplX9Vt8N2CaY7HzmrZyq7qDqWxc7L9mnGAqzOH/IAWAYiHTttMWzRiMyT/7EYt5z3csVv8eU05P0BtJn6XWHE3uGnpYpmJbPdGysaavhc3ZrPOP
Lbo+Vd5nJ7VfCfIbjwSwZ+g81KzuoYdrw540abZft84VhlD12jegMWWZ8SIN/sb9dX5paOQs+KvOzMXnmng+vpcVCcpn6ezB3Fi3lnU+qIBL8pfo7E6YLfUEOgcuPvM9
pChKrE/CecFd53QtLeicr1GzKDTeWc3lY/tIHJjNxgwe8Ov7fqfXcidZmkSpqikYyGRI3eEO+6w7YLsAvQZ/9qPChihdOOnpCwONSvvnwK6BEqKLIQkH0alApiLWW2Il
j/lllaamehG399QiykV8HfLWESjonfi0urb6sPousqs3N4SiLFFulNap0WZJ9IOMwFghpdL6dlJbdeuePkXrzST9rhK86YmwyB993b3hn8Peq25dQWQGiK+Q9CGQ1niB
1m5UtOi7EoPtaB+okLeIHRlwodcbVYeoAMOa4jJzf9d3nJzPAwJsYU/ZFeUdfXGSOwrLUQIm8jVzma/03GBkDf2AK3VvBVUCB3ltKEI2RAjIHJqn6UQnCR7A0Mq17RZ4
2OPOJ8nu4vgs0Z/doirk8BMTJq6vKSrtRmZdASEmvZvabX/la6jNG/qib09aNdKQB8lRZBoeBsWZiTO6bLjcMkvEcR9DuBot5ywixm8p70P2K7wKz4HQv7ab6BksZNVC
/3vQwyp8Mit6vANbO1OFpj0kbJnL3Y8eQBC7IV21Ef0hSFLTJJ1RD0DoWVeb+JFuWuQwXDv8+EdeRJz+eF0ZD8C/2P5yyD7PEakQ8tbcaQZ03g+SrgioieyX1t78eFyu
zmhHYjYrWLLO5EHpZPREXtCVzrgH4wVT2nFuXRdGdDDURmYUPjRqNehFAOUhvM7mkIZ9WFEEZM3tlCCfWLs1KYv8J8awLNHuiHygEs1n/595GM01SxMwHgE5cO/PDztE
FI5BmP3nQmitzDDoRZmdvq+ggEAdZ9VDtPNDrreJVZrnc7HGMu5kB7sM8Mx0JK1Vx+KTHrDWLuW+pwFHtNIi9QfJUWQaHgbFmYkzumy43DJLxHEfQ7gaLecsIsZvKe9D
7fiKNaN8SAs3CvrMR59hFp94m869WG5dZDyjdD4bPk8lRw9iFJeqaWyZrceZPhk7ZIlOTpxjqXliYsYaSvUraog2KG8sG21WSnAybqd90zqDt63YRQAJMndOEYBkjevb
Mt7oqvQw8yKBJPqR4GgQMFhczYY5SV4cfw9i2Ac6UPXaFQ0QonvmMW1hI9FBO3L6Ump0qAjT7YgX9v1rw7WqJUQmqywOJT/O1QDN5JTHKliuy2dKbe/laBAIN0D/6LuB
5+oYCaTNVp2vZGkvMggUWVUQEhoK217dO6xwx3++2wmRybAyhKjM97OQqLMXA00Eyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iq
xpnyhlTUUhknz/XpDdrosB5y3ONtEX6heqMlYyFdjkDKiCbRJr2HgYyrX3ljAm2I1Lq9siTdjb8DHmpPMkhZYlTGlDJ3QcBfpMDJLF74XkbKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiAYWk2wHbar4ls6j++L3VLEzPPzHWtnf3OQhSyRuWEvPoH0QvhzQYIzWdu45fQ9em1bqzTfydZ1dAcSrI7PddMqRUJgmvoSRx4YxQ1jt9X8V
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L309D7us/dNj4/k5+TojwBuHLt0O68I/LSrTXFVnixB7KiCbRJr2HgYyrX3ljAm2I
bAeeCRycsmvOpBE3PLXopcqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IcgcuqXz8VKFxDjVJUfNjdtyEK9mErwTA6gB+eOSxUjJOhNqhIcdXPGMrmn23d9Eg
yogm0Sa9h4GMq195YwJtiP72e5pQo6xSGF/ma7NAvnnWimvusHDbyMQ41+dZJGiaUOF2rAbDcUn7kJfZRNs/NsqIJtEmvYeBjKtfeWMCbYh34VQFdncvc4rGqHSJ35gM
MUG142jgE2cA2lJvjcf3AFMaEHlsnQsQyKZVFILUEq+CymdKNs4MPDwvtFZYfXzupxfc7XrnmrT2eWXhTEq3rMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
oFN7gHeT+ZseMhR+qjrtIvkt6AndwIj3YkE/k6qfXXoFF0ppmdU9L5RUDz4ApzFpyogm0Sa9h4GMq195YwJtiMy6abn8/DWptZueN5oEPKgZPW5YbP11+pb9eGjIUjZ5
yogm0Sa9h4GMq195YwJtiE9AHUqNPiKMXd6TmqYHnDFClrpE2BmSvu8RxVfeL5Un2CBNR7ngbP91VZ+4oskCoE1/dFQI+bNoTdA3CtXKYvTsm6QgG+Evpo2JgZJM0q28
+1cAfEsrtMMr/DjKV32HTpDzX8clJ0r/8Os5RC63gPfKiCbRJr2HgYyrX3ljAm2I0vZ/C5D4uxV8hGR06yAxc6u9D0u7Bu9sOwgU11Cm/95MAmZrmH7lBkJmHmYs2DNK
Ko9m9Kwl+fV9EHP8S9v7itgkwfW+J1lI+OHKXxBfogKYf/OiukdUyTHrIJx5maW6yogm0Sa9h4GMq195YwJtiDZlloNdhddpYOAaTVdVPMefq8R6Aa2HFjgvab4xw9u3
7sx5oLVAd7tGDiIrzv9a7MqIJtEmvYeBjKtfeWMCbYgSUykWX6EgCQ7U6wPFhr54VMaUMndBwF+kwMksXvheRsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
BhaTbAdtqviWzqP74vdUsXHzghdMIbJedTNKiWQq/xkM13OT5sTrd78r8JRwGuC2YtodNI6/BE/oMLHVVoKgQBuVCKJu2x6+BY2vDbvErZ8odpT2S9d1sN1aI2EbuFh5
SQzJmoDESQr874F9tLs60YmvX5jRYBoyP+S0/fQvdRrzMl6y/FwkogN6Qi5rLRO5t1p0CWaZhrfk/DR5adN2CMBlLkdb/0BuAiSXEClshzPtceNbkK1Vtf2NYkzMpHeQ
rqQPIMZHQqeI1JCudQ4FYuilxajILmjYeo3tjVwCwlU4cznkjkYgROsFqXIzY+l9PBKPPeV0OFQvvd8o8dKTZqKUiIALyV48nDLVES7GDhZpqBKEqfEf6cDmCtWyUoa2
WU1HIK49eIz3DYTqG2kQP7o66APqRMr+xVZjnPk/m8YJf+zJtiax8l75189ZOznxso/gQHQzNSGgI4dnl9eXdca1omAuN7tugAFrz+M154t5Bqj2VnrnXf97uo/5DCdU
awwXqJIiEQ2Z+cTdiPERWgXKksjmMPHyKFg+j404PcM3l8ucY5RtLl1XIYPv588WD5C8fVp/xNbB/Mxx/Z/bI7+BWpAakSEhauuNrRlVl1CgU3uAd5P5mx4yFH6qOu0i
+S3oCd3AiPdiQT+Tqp9dek74DJrsd0fMjuaOom4W3jGrJQT6sMDyhGAZdv4Bjxt+I/MMohbMNmtxkhXKBgQ/EcqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
T0AdSo0+Ioxd3pOapgecMUKWukTYGZK+7xHFV94vlSdd6r4sepZIAksLTH05b0GwNyspp5Rs+l7Bbbqs3gAxLlfW2O1xZro3ekCdoofI5Uf2d22BCzSZkAkBGWlH5aTE
yKjVqoO8cNQWMkCEm+UqJcqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFzhsUCmqmG5eSSg/78P43u+zidkfumdyUkifGYwozI852YGmhumGUMxdjMyyVOV2qp
1opr7rBw28jEONfnWSRomm0MBrnUZ9YY46T2wBcXz75MAmZrmH7lBkJmHmYs2DNK9eAhsbYpcvuVPp86ImPIqp+rxHoBrYcWOC9pvjHD27ek3NAUIv2LWDGDnjNczDrt
9ZHbzlBOhOFMRiwePwts1G6zzV7+LIe0z8muPQV59OuUQakWoxTwHXjA1UVKJvNPXOksEUDfNp1+QxwTX2q8LcqIJtEmvYeBjKtfeWMCbYgGFpNsB22q+JbOo/vi91Sx
cfOCF0whsl51M0qJZCr/GYid8NDgNmWWWT5FtYUNQWXshbpBgCjk9OW+Z73uG5gzDbYsu7C9SF70UGqlhG7LBQghvRHv7F8IJqdiM7MQAa/KiCbRJr2HgYyrX3ljAm2I
KbAWmvuvd8ilV1icDV9dy/MyXrL8XCSiA3pCLmstE7m0Gy3MkKs03TlVupRSr/3txs+RNso6leQF2yCntJEJxbMoVg/m3vTC6t7uwKpO/xdY1SzqQ9FUzVoz8kOF7sE8
I3gCwP/oPguCZTLfoPZ1DnIHLql8/FShcQ41SVHzY3bisN/Sh2n8mqpk2ZpVWHHJpv6cyBh22ge2q/yRPqxLEMqIJtEmvYeBjKtfeWMCbYhCIOdhNafeW1u8GGt0l8U7
ujroA+pEyv7FVmOc+T+bxuzx43Af+A9Ds++SWVapkBXKiCbRJr2HgYyrX3ljAm2IxrWiYC43u26AAWvP4zXni3kGqPZWeudd/3u6j/kMJ1RFOL7yaxmymVIO1V21MOUO
AivsW+pKty1L5A7AdtAkPTeXy5xjlG0uXVchg+/nzxbcYM7sLSCAcGK4AHXmh5Jdyogm0Sa9h4GMq195YwJtiKBTe4B3k/mbHjIUfqo67SJIIXCDXnvXctbZSEYRJJYF
Tof61BeuWfqJVRDNP1+GlMqIJtEmvYeBjKtfeWMCbYik24FGdWl+bb0+yv3Yedzoyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhPQB1KjT4ijF3ek5qmB5wx
Qpa6RNgZkr7vEcVX3i+VJ5+ahOjsWaN+fsicNaSljkLMEOrDFGST6DOvm+tIGKSJ3mAFi312V17kTOEx3HqBvikZpRaEo2S3NbNhztSaGwb7xGAHupGIPjCoXvFZ5ObW
yogm0Sa9h4GMq195YwJtiNL2fwuQ+LsVfIRkdOsgMXN3EkF6bXf/Q1hQ/3NbSvcizenqmUNQZ/7Fp9Hu/fQjuFUQEhoK217dO6xwx3++2wlQnEMthiv5vDqFF/MjGnqg
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iqYNbsIYA/55OXPv6bZCUsU6uIDGdz+39V+KuYdjkqlLbKiCbRJr2HgYyrX3ljAm2I
/le6S8roDXvUQFOq4e1XE1Ok30DyyuJ68QZZntWVAOQog3wX7Md6FpnuFkJExBytyogm0Sa9h4GMq195YwJtiKvdJGLF4X6YkZZhiH97F0QlfR9fxmJZOtjf9xh7/fFE
3MH3yNHRPOMmuAV3JC21M2LaHTSOvwRP6DCx1VaCoECGl/qLjFuUuh11A/9NIeGyC4/Mq49wfYeC8zqaroEUDMqIJtEmvYeBjKtfeWMCbYiJr1+Y0WAaMj/ktP30L3Ua
6a9fu8vaeFkVZ3pXoqGYyc2NyfjyLNSnZQyigu9t5cnKiCbRJr2HgYyrX3ljAm2I7XHjW5CtVbX9jWJMzKR3kKp1sygJUJQ3Tv+H0WLNLEVK5GAQ9xk1ZRdGxNbFTdoZ
cgcuqXz8VKFxDjVJUfNjdgittQ5KvqJo7QWFThbpgtKzoB5vUBuY5aIzjKAIElkpyogm0Sa9h4GMq195YwJtiEeljPCPfEdjrzZyvRwc8TVjiyjfzVTPXrFbZ99I+uLJ
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYh34VQFdncvc4rGqHSJ35gMzFqkkAIUJ49NeA7vfOdOH2AThRtkILDS/T+x0zDWjrLz4Z2jts2hgE3HNoJzrtrx
NqpSj8ue9wBTnXr2BJnmPgFFPY3B76rtIGQEkanXBEFm2MOx20XdI6mdxqOZ5b1b6cdV+3ONhDnp7Kb9AzvcQkghcINee9dy1tlIRhEklgWjTF6+dnaWnAFj+HrYMxrf
OoWc0EFu8wIwBcC/YD6kzqqJZW+9tM7zX1Wiji2GJ+k1191b0jbD9Vi90/0jHXWq6esKQTCI0/NUDdcRkl0dgk9AHUqNPiKMXd6TmqYHnDHqDL/ryjNec8xTlJz9d5ov
b0RGe5bljJkNTfz8XLOdUxkuM1fh2wv8kMnQup1PixTDI4YLLvc+Ir2GCDX6YxvbK9CzmFe/IxyZV/Qltvwax7SolByl+r8fvNRgshaHl3uBtdaRBqeOTD5UUzy+4K+A
ql1NB7U/njFU5faCQY2X1ysShiFGFUQK4eZM0TyyzSfKiCbRJr2HgYyrX3ljAm2IKo9m9Kwl+fV9EHP8S9v7itgkwfW+J1lI+OHKXxBfogK0vhLmntq2hozFZUzsuAyW
yogm0Sa9h4GMq195YwJtiDZlloNdhddpYOAaTVdVPMfCc00dp/uVICRuyrwaf30MT2bdAfGwY8ZDwAKPJZG4w8qIJtEmvYeBjKtfeWMCbYin+TQ7VCrXq/F/EfaUItAy
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2IBhaTbAdtqviWzqP74vdUsXWUvMeKYXArztNDFAJuW1XKiCbRJr2HgYyrX3ljAm2I
YtodNI6/BE/oMLHVVoKgQBNM7jsKa69JUY3Ni+y72ufj+PkMZgKZDmvR7ccXURbDyogm0Sa9h4GMq195YwJtiImvX5jRYBoyP+S0/fQvdRpOq05RAsAcjIXmWiy5LFEh
yogm0Sa9h4GMq195YwJtiGfhCgebeW7GZjswfY7sgyYnycArXlCYlBQeiHAsCVvw88JKhJEpeOwRxLuj4ic/RcqIJtEmvYeBjKtfeWMCbYiJr1+Y0WAaMj/ktP30L3Ua
nD0420jKJWnjZcReg/SLb8qIJtEmvYeBjKtfeWMCbYhS05M7s90EhofheSI9h88awPJ/mWDwlvSlcXFJ3jyJdMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
nkPELMSQBI3KYVRngPExRnOUcCC3F3Z7CvsLtFXLw+rKiCbRJr2HgYyrX3ljAm2IwyOGCy73PiK9hgg1+mMb2yptcfPCnfQSkX+5icEaftLKiCbRJr2HgYyrX3ljAm2I
oY4ZFtMWUeI69RCmMkyCzUxSaKeImIhfMmL4Q616D5BB4HrjsQ3G5b4zaNKkE2VSwyOGCy73PiK9hgg1+mMb2zpMrZSYiPQLyBGX+faaKuLfQMlhF9m/0TbE4QWWS7P1
oY4ZFtMWUeI69RCmMkyCzWbEOeuAgmsa6wwBRxLX8ERShI95T9PkBrwcFddpZV9YwyOGCy73PiK9hgg1+mMb27TTFAKv7XFEOPau3nMIl+DCTAURt69yux/rAUYscbHi
oY4ZFtMWUeI69RCmMkyCzassMPCmTlPoDzCo2rQMNnOIk82ngUM3c9mxfKXeXDQywyOGCy73PiK9hgg1+mMb24gCYtoQrQs1FUOCnPnR+gAlscb5OtKF6LsbG7Plj3im
oY4ZFtMWUeI69RCmMkyCzVJA694D+TAajQsQklGFpymKHIV2tXiGesBOoq7R1Q1ZwyOGCy73PiK9hgg1+mMb28qJQnH4/SSoCFQmD9n21x9giNjqEPAiw/CoQUIU+0Nd
oY4ZFtMWUeI69RCmMkyCzaT4SzYfgopLlv5pqFfKT8YuYpGIjaUi7tf3s84xauPrwyOGCy73PiK9hgg1+mMb20n5YCMaFN8C39EcRvzNOkwuYpGIjaUi7tf3s84xauPr
oY4ZFtMWUeI69RCmMkyCzTnAQhzqvW9TnvyQ/goGeYn7rICpy6vrQuFpgCGDT3b1yogm0Sa9h4GMq195YwJtiD88GAsZtuxeUqq3wSLdfQL6J5L7yLtUx2v0JcgPkKuY
yogm0Sa9h4GMq195YwJtiHIHLql8/FShcQ41SVHzY3ZbXy3X5pc+zbiBjjbnx4gxCo7KGgrEloYK3ibIw1o1kv+6TfeHc6CWg6mFbIWNgY5TKYoI3sUQrWU6aqT8UpSU
uSPfxyv7eccgSfgeHT+HJcqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOejWsk7MLeHe4yUrbRfg7QjlsqIJtEmvYeBjKtfeWMCbYhvRkkikjWh+NVzgLgaebmY
6fwWPsY1p4AbJi475Le097L5Tu3BJ0g7sMZt1RohSNfKiCbRJr2HgYyrX3ljAm2IhHN5hH9F82XlRyJS8p4fpUwAmsMeYpW4YWfGoZsD/WnKiCbRJr2HgYyrX3ljAm2I
YNLYKxdBjjxtb6GvKOUTFIiTzaeBQzdz2bF8pd5cNDLKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiKoGj5MN2FrbDQGGH6xddEs3c5wuSWL0U3fW+ed3JyVW
e66gG7Gq8vHYAlsRz9zM6YaOAZNwhn7TueSbY4xgpoDKiCbRJr2HgYyrX3ljAm2IQiH+6sC7fVPv/ZRtl9Kr44bHHev+nNLDPb+xB1nQJpR83UNojvRdbs9N03+sexEj
NXHZLiu+/k1w6ZZ7QcLWDYPIpPUGGzqUpTZmAHT3Udmn49LTX5XyGNoN71UBz3U/yogm0Sa9h4GMq195YwJtiOyklcPwIR6cplmr8SC13d22+h8T/WUi7sjW2VYwSgEI
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjeBEehDRu5tBQw9W4ARUw6Rmr0aVpt92Hr0sNfT6VRH0/r/LY8Jexi4fmcI4d7szf7rICpy6vrQuFpgCGDT3b1
i7nfm6WPfYAI3VWI2zNP4cqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiE9AHUqNPiKMXd6TmqYHnDFClrpE2BmSvu8RxVfeL5Un
knkQy3asTOLRUghRLkcWzsqIJtEmvYeBjKtfeWMCbYhJYxC/pojLErGLqKPmZtF4WG3e8Fuq5mXP/aN5hHQAbMvevs6j1bZdg5Mwz7uzgEqJCmlErDSoIVMtKPsuI4yD
0yGRnPZE1s62DA8g752IHMap2fYsbBVw/U0AI2/Wuct70OIh8oUXcyDJ2flr4ZqHyogm0Sa9h4GMq195YwJtiJkqZfjZiNJWu5Oo5FVmDLlUHx7Yr21vdfI1oZsZYkIJ
AeuSDD2BdzczNrTXqwLwWV48xzwfEbNlxvwSufHfiKVyBy6pfPxUoXEONUlR82N2jQO6poVr2LWu+Tsii3hAulWouATPRjWqLASK7WKbnEDKiCbRJr2HgYyrX3ljAm2I
0dzKF/wYiRK9AOq2Y83egcqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiINxF05+fMMIhjTy+zEu7XsX+ojaUT0RybKFhISy/4pO
WaeAygVbvjPazzznEZISKcqIJtEmvYeBjKtfeWMCbYjTLUGbT+kdmy92Qrz/3GkByogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
9eAhsbYpcvuVPp86ImPIqqelt/+vGiKltxuYPdccLfMsYgVBpvWw9/RauHwPAluEyogm0Sa9h4GMq195YwJtiD9q/bTkuFKxWr1Vsm3NH0Fz2N1gFJXKiw86AD8xAKwY
OP8FoDq0i1xV19PKzLcyqcqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFGyR7BBEqeXgyxZWuEdN4MU5EmOLiGake6w3XuQS4a9kHKiCbRJr2HgYyrX3ljAm2I
VTLZGq1ok0CTSdQuWGlkQbwjCYbR4iNwqXDZa6KRsdqCqEw8b5Dhr+5TW5NEU6eb9XS9Exuf8d4wnALr88gMnqBTe4B3k/mbHjIUfqo67SIaMTkhbXWpuzysYdAoSAgu
8FpnaOU8oOxbgtDgG8ilO8qIJtEmvYeBjKtfeWMCbYhXfU3DausIxILYlQpuW5sspA5rlaC1sFOTZ6DPVgB2svpFw+nDnnGSX5oMWUozIr/KiCbRJr2HgYyrX3ljAm2I
fUgoSjZJ0mfLOvTfraoVzuL5+35c1RBh826gyj7+Cct0RSA+lPHlnGgJunDyrzvK+6yAqcur60LhaYAhg0929aKhJvYvdC2BgUCoDMBq0RmvGtowI86xDBoS6/L7mZUE
2gHGDyxsNQu3F7d+hAO180kMyZqAxEkK/O+BfbS7OtGJr1+Y0WAaMj/ktP30L3Ua9UqzRW68RNlOqoAdoNq8oRmSjCqP1bIwHZS3WF53MwwPmZNq2ClMOQAHWKCi9Jwr
JryprLDsfWvjd9IOaMsRqKiWUN9fztCslafF/aWbqs/0SL05cIzYf9d0CJiGiGQF7UVSAI93dHdekXcCTfP6gJcxlX9YO+c3TxxC0LDHZG6BwkmKaj4tMf0l/my/+CEG
6Db2f8tJjC+bTbp6Az7iTOSDtX0O58hQd4tbjLy7MufWimvusHDbyMQ41+dZJGiaVrgUVDeYlOTrTmp2oFGOCicJZPharvd3HVwikwBpxsi2bEHb1zjdym6SuXY+nEm6
ql1NB7U/njFU5faCQY2X1zF8Sjf9nEZuCn4GSov0ndYUCgxGjtpU6X0c10//kfJGCZxGhU9fdMOpx43vr2Df2ir/pysRRcgK+nqG1OAZUmdkTkrrb1WX22J82g0uyBAN
x9rSvFJKQKJlxdCXLTEZQ8qIJtEmvYeBjKtfeWMCbYhQVwys3bC5W1JiegIIlSi8EDFLetJXOtUzBdiKqkHViZbBybm5cmI2XNvzl9KFJUR7O/cE3BUYGSGN1+jeXx2+
N5fLnGOUbS5dVyGD7+fPFrVsh5SBjr22Ws1Dv6/MoGeJW6BeCc/5yLB1TnoGzvIdyogm0Sa9h4GMq195YwJtiHfhVAV2dy9zisaodInfmAy1ynztqSgsSgYLpFm64Chk
ivfpMAL7c8fjqJg4l/1FyREkvF/ruXc6VY+hatebM7+bHyT9yFWz97OSOS2+RGqy+Kr3Kt15vwPY8z5qsFaTFE1/dFQI+bNoTdA3CtXKYvTKiCbRJr2HgYyrX3ljAm2I
OmcBZVUeK8oNMHDzLDhywctNMSB4CV1fcoIEsMntlNgNyjBWVPsGNrhEOBoEg1d/PYr9omQjyb08DUN6lnUU/Q22LLuwvUhe9FBqpYRuywUwQBZ/5kq8uz6CYO4ecIr1
3tg36JZIjTN8D7VQ9R/VssqIJtEmvYeBjKtfeWMCbYgGFpNsB22q+JbOo/vi91SxgYpdTorC6Lpc9i+HPShBL59d6WUsxYoTczns/5gu1iWaJvXGscLNvgOZgzQB3C9X
X7aLw9jhUcNJ61wZcmMaWf1aBFdddMc6+dPX3cq1cjF4JiCj9Op3wSb5MCvg3JO63gRHoQ0bubQUMPVuAEVMOkZq9Glabfdh69LDX0+lUR8AeiQwuQ3ooFfhg2F9TTKo
G3EROU7t6Umug5Z7yeVALaFrHFFSaau6JdAhGtmzznf2d22BCzSZkAkBGWlH5aTEiJ3w0OA2ZZZZPkW1hQ1BZcqIJtEmvYeBjKtfeWMCbYhPQB1KjT4ijF3ek5qmB5wx
Qpa6RNgZkr7vEcVX3i+VJ5z0ugnL8/AEdgZY+zcRSydp+3F0ysKd8wZbJC8CYnFsSWMQv6aIyxKxi6ij5mbReLm9FA2dKk0jkhVl7Lapp7TGT/ZIXMu6w3fGfmwFvzOg
yogm0Sa9h4GMq195YwJtiNMhkZz2RNbOtgwPIO+diBwNvhmJFnden904K0T9vZyraiLpmATzUUsTLC5H7N35ucqIJtEmvYeBjKtfeWMCbYiZKmX42YjSVruTqORVZgy5
VbcC6Tn8V24xFIMZ8VT/GbXKfO2pKCxKBgukWbrgKGShUTnC8uHvZX8SRiJq4JZWcgcuqXz8VKFxDjVJUfNjdqhqttuSRRKxX1HgOdNw2jXxFMJHWZp61KR/cMzjy4Bg
yogm0Sa9h4GMq195YwJtiOiXtY2LEotFWJ05dHCfwJzc0Prq+o7ZgLrwv/mT9c/dYxlBvQct9YC/FcUwgojRN8qIJtEmvYeBjKtfeWMCbYiDcRdOfnzDCIY08vsxLu17
F/qI2lE9EcmyhYSEsv+KTtYCV+scTPHdgOvImLnXrsCJW6BeCc/5yLB1TnoGzvId5CTSeMLqHobmYe6Y1kpeOxusdyBQHriUPhu/8nLxUViUiSCxmGSdY5Che4UlV286
v4FakBqRISFq642tGVWXUDZlloNdhddpYOAaTVdVPMenpbf/rxoipbcbmD3XHC3zv52rBrPJ7YmFwfRqAAcfpcqIJtEmvYeBjKtfeWMCbYg/av205LhSsVq9VbJtzR9B
iczLUsL7icy5m16oG5CbUOR9LEiwEoMFM5EbksbQ6xDKiCbRJr2HgYyrX3ljAm2IoY4ZFtMWUeI69RCmMkyCzVMYZrPTSc2pgTpBkXeYIql9bPAjTIJ+PeKJysyrv6lJ
yogm0Sa9h4GMq195YwJtiP1lXM6BWafEAcFZCxPlhX/KiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYigU3uAd5P5mx4yFH6qOu0i
VQacVG6Mc9nsEOUTQ6Murbtu6PFbdvhzOcW3wsyUEhXKiCbRJr2HgYyrX3ljAm2IF2y2DBs/HYxIeXpe+kgedMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiIEayJwYGQ9fRzfY+QWc56OA7ZXaGw1oF7JExFujDK+UBUDVp+gfGVd7h8jz3x2+CsqIJtEmvYeBjKtfeWMCbYiioSb2L3QtgYFAqAzAatEZ
E2jAl2KbqYJcHYVkWCpkdjHdW+BerXtFaJHnc7+6exO90MQTff9j+jv39BdzMv9pKbAWmvuvd8ilV1icDV9dy3weUbw3LYCjfKiVNkjWz9yApWXnFdl1Kf6dAufmT1gD
SZXdRwN4saED/s81w/rdTCa8qayw7H1r43fSDmjLEaieOZ214n2/1iJeXx3IgEScSWOBzhjuM87v78x251kze99AyWEX2b/RNsThBZZLs/VAyaqwkAgzq4ApJkwTRqQM
s/laDAoXuP+jd4jlLJEkCJRU3KrYBA8P2S8kHgmM6yno2ACt66DzP1S77w/VpsQE1opr7rBw28jEONfnWSRomtwUwtrWbhrBNBKdS223buDdSrYNwxYLBtRem8MTDxtq
yogm0Sa9h4GMq195YwJtiKpdTQe1P54xVOX2gkGNl9dVIDLdUZjy8jqmou3wZuQbqo5PHIm3vEF3VWugaLS7JC5HhTylSQQAbQFVoMdpU9E1cdkuK77+TXDplntBwtYN
H4MqwX9AoBOZF1bED9lbk8ddkRW8MvgNkTcbASXN1iTKiCbRJr2HgYyrX3ljAm2IpVd3zd04KWktD7F0hC+RxhWURkSy9fBHGc0HyKvrb3dg/xDfzwWfPwKUImh2PgKK
wDttir92jWfwspbheHTF4PzF9rwufWaZBQOGyMy0CdXjasVVEM3aDlcLZZcR8iol0NG1+UEXxH1i2W5u73t/18qIJtEmvYeBjKtfeWMCbYjGtaJgLje7boABa8/jNeeL
DWsSNq3YyFcIS9avnyTQk/p1OdoAit2U3WiuGRtqV/ARJLxf67l3OlWPoWrXmzO/TNRs9sZQQ8JaSXBa3ar4MQHp7t1OxKQIWyXNyuwsFJc+zuTMnVyznL42Nx+8rUqI
yogm0Sa9h4GMq195YwJtiIUc5zAXPCFOpd5czvGFIhQuHOBh3YQb5A8ZGimpIbIJiKef8Le8NW32/DbaTVoADT2K/aJkI8m9PA1DepZ1FP2H03VxIlv8vDyOeM3Rgw64
lBAKB64FjgxYA1ATyHPnzJjYz9HEoh6oFQUD5W3SuTjKiCbRJr2HgYyrX3ljAm2Iq90kYsXhfpiRlmGIf3sXRGcJlZq4ORojRdDk+y/JxCTKiCbRJr2HgYyrX3ljAm2I
7KSVw/AhHpymWavxILXd3Wx48pws7qHHjLkatVbLFoLKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiN4ER6ENG7m0FDD1bgBFTDpGavRpWm33YevSw19PpVEf
XIGytOXTm2Xiw6I0Zq+oLcqIJtEmvYeBjKtfeWMCbYgcxjFVBlKGgARYFh2hxll0yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
T0AdSo0+Ioxd3pOapgecMUKWukTYGZK+7xHFV94vlSfLmZNmMXKqd+8lpreB/Jjxyogm0Sa9h4GMq195YwJtiEljEL+miMsSsYuoo+Zm0XhYbd7wW6rmZc/9o3mEdABs
46DS8+wVKqt27Hknj2Yrga/MunTTRkY6ABEOxE0PKWQnHskfB9QusOl2qjoY4Mx2XeLwcuuIJ0aoFLzhxwr3v9p8KaxIxCfwRJJPZaJ4EinKiCbRJr2HgYyrX3ljAm2I
mSpl+NmI0la7k6jkVWYMufE5LE+Zggq1pvoNvgTC6rTOgNn+h0jGzwupwl3UCMEpyogm0Sa9h4GMq195YwJtiHIHLql8/FShcQ41SVHzY3YPnKXwm/CFJ8ce3p9cCQy3
cO9FJ9UPSFHOhvdRrHl1wMqIJtEmvYeBjKtfeWMCbYjfM9RKufRLOQSEDQb3VE0HcjveAzO+/7U58YwS7JUaF8qIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
g3EXTn58wwiGNPL7MS7te1znkec08mZzjkH4p8YaMpH9lgUOgHfDiJgif2hoMD+dyogm0Sa9h4GMq195YwJtiOQk0njC6h6G5mHumNZKXjs3Xu/P+Eum8KWl8Xe5CH7c
TUbcATlRf7DVWvJAxKswkG49yqOPgox/MoPbrhsZmZ02ZZaDXYXXaWDgGk1XVTzHEeJ4i2Y2jizO0/6P5Nb1Xp6baVfWFnCoM0S94XgfnyHKiCbRJr2HgYyrX3ljAm2I
P2r9tOS4UrFavVWybc0fQdOYSVnkHhPmyWXkm3MKWjOKsZjxspRdPlvfgkygQGhgyogm0Sa9h4GMq195YwJtiKGOGRbTFlHiOvUQpjJMgs05wEIc6r1vU578kP4KBnmJ
+6yAqcur60LhaYAhg0929cqIJtEmvYeBjKtfeWMCbYjsMQIHiyCIWwfiaOSNB2mWTX90VAj5s2hN0DcK1cpi9MqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
oFN7gHeT+ZseMhR+qjrtIp4AfWdITcAsp1PAuzH9ySTKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiC/Nsw6V7tBXW7MGU9j17xKWYnCpLHNzGAC4XS62ftEe
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOejWsk7MLeHe4yUrbRfg7QjlsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
ORHjSbjCtTM1MGQfHmRkZsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiCmwFpr7r3fIpVdYnA1fXctMnmBDOkr+MD/K7wAq2YFr
yogm0Sa9h4GMq195YwJtiEmV3UcDeLGhA/7PNcP63UyAZY1tUInPvwM61cJnATUByogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
9rswH5Rl3UkeJz+f63rT77iG6Hh7LEqB5xE3OGqv2X/KiCbRJr2HgYyrX3ljAm2I6NgAreug8z9Uu+8P1abEBNaKa+6wcNvIxDjX51kkaJq111WOJJg9JuUFqtHnlfwF
Vfp0FV8VrcqWlrn9wo8DXcqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFzPvUdOfXibzV9DL88htA2RMqIJtEmvYeBjKtfeWMCbYj7GF3hkVzKZAoM5pJGg1Hv
TACawx5ilbhhZ8ahmwP9acqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiJ0Wl9N2kOxJrtSzwsuUoTwhI2xI0PItUgvKKCeHUfYz
yogm0Sa9h4GMq195YwJtiFDadW6ph1b8t9G2UQNc9v+Ao79L2BhBoQd4X80WK8R1yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
Mj+7Ig9yyIKuNSVxrFsJmidS0pxUvTLXrrHlBjMFDCuSkurkf8fI97kWxUpCAw1yzgGacj1HHzCR5yyJOstzmpuzlKcqq/ao33z3tuzsegJ1Pa6XoQ/nmTRn0qHRCuhh
1opr7rBw28jEONfnWSRomtJ2VoR1tCCKFkeo8eHAVYeQJ6umH5HvmbqX9mdtaVSHt3+eq9qpknE5Kp4VpkCCbFzzsg5NyAtJpOhm36VgeNS075bSc4EkOT4TCaRM5nDi
9CGPHa4mYd2DJFbC08MsbPrxGf3wSKzJ1Z1GfcY9qHD3rUqOOiTSIdhTIMg5HViu/mSQT98RqK1NHuNV2iI7Tc3bNu0gJLss+nJjcYhLwlcCq6fhhj4ofux1kS1MBH3+
GTq9BqcEqrSCqweEMHGM7WXukv0HH+aCk4I9JrjGZAFsOdeMw+I51HrmG1xMWvKo8p2FBN7SzPVTGIYvNT+7ZuvbSK2PRCqHBfn/CUSidOSt4U1PJ1eRKmyGCSG6sfIz
GMFu48Bu/TQL1ILJy2CuJiaB1vvLZumnli3hXfK+F784QghyoTFHanxF43WbEuDvfvlpS+vpSmNu4ld+HTVI7zv0PKof5FICRQOyETz2+vMwJoq3eHhJnelKsER8QXpk
7gZ06FzFmc39GdQEc7a80u3A0H5QMHpF/iW9gcBUqNFrKEs/b/4ucsUKwNuS5Am3amGMtAQefMD6NKK8AFhRtcVVXUZyh7BAHXM4FoYUCCjOvcruHQFeZM30kr2GULpY
isX56zkqmBN2xsqiy3C111OnJA07YfjZZOaFA29WCWk3ie7WOvFaIFNMn/k6g8OJv9hVj6vUGEkWxB0GY5HzYzCtVkgq5Yl9Zphx+XBAO4kGV8lwCa0/ojbjcb8lYJ2H
6GaQ3Oa5vzb3oDM0v2yB/9rTMApUhmfq6ZoHS3n0yanaaGNdww4Zrix3EuqQDoGnc5fJFL9VzLZIbD6h9BnvGAbfJn9hWCz6jOYXszGbmq6b9YMzCZENTTuJ/skiUn2I
M/sZIiHxz+T3h+ni+TpQIBeM66sJCjBqGBFAK81OfKjQBfDa0GjQFlitK6olx0tmcGMAqdfAvYNdnpCn2ncawrniZSs2iCi7ZeesRoIQJFTQcgmCNHEIqmlzBTnMdMjR
ll0dnW+rsp1GahedloHVhyl2/IqSo2Dv01Ko4dFJwZ04z1TIqVcHQFIYFQs5cOK5auX47fj4t6fqSnJb9VuZ46YH7C802CkdXmOyVN7y42ShCTvjSxfmlZW/LNgICIbL
QNiFsbz2gaTpWeYGTFAF8V52C2tZbiHmsMVVnA80zXzPPrGR47bK9pVeOQru7FI0Y4Xs8Oh2mcce3aa8nbmaem4T4kfojaO7PkeslMy4PcCzmJCNhcuf4t3U0zKUpCqX
qo/YFf/VWk1d1sa+HeHpCtkx/niARTtdOrk2kuko2nE1gLqX8WBS3xlzRMp3wED2J1LSnFS9MteuseUGMwUMK/vDtfZiMvIaBM7UAPhQooqoAgCTEZfQD4c+SG28hCT1
pQmXGeyj/QjmsZzaFLEmsA8HwhdfpX+cNdFPLgfrfQOWHiuSdsLWJRyoVM2iQClFPymQWP3awkMPYvyM+oN3tPn+t/cixky4oJxmx+gIPN+lCZcZ7KP9COaxnNoUsSaw
dScwlH8lf73nZMV5a4MhFUm0GAzLou1j6Qcrb/14qYU7+MQhZ9kHUQAPofMsku09EXfLgORrlF0cfLvRwwV/Gm9kTp9VOLwMmhO4KWv59SfV/mC2/O9u9p0uXHicJ5+c
7cFPk4BidCbOPJtmB6UUBLF81t5lL2YB+PoapISPPPfh/EuKzIy47gsKqbCnOgtdBt8mf2FYLPqM5hezMZuarpv1gzMJkQ1NO4n+ySJSfYg3foUvkwKf1K5eGjc5Ae+l
ysMsicYMYkMRgOD9wpv2dtmHfZ1x7NfUPlI97ivKn87R+v1aPvQfZNBryfGaExkvln9Xo+sW30+qkYHiTC2CALOYkI2Fy5/i3dTTMpSkKpeF3tInMl5eUr87puv8Z11n
hqNGQQzqgZFA4xsXg5PcEV24s/tScbe3QG2umSXFZPN1541jkYoAbWqKoJQJmX3o4P65Qc/yIJWKGyi1RxB1bnR0gdvHwyyPygt60MLL6hwi/7jOWDh20YrHw+4AuYTy
yizTFVTkFPiJ+ZAsu8F2B3Y/p0WxjQv7/psoxY8fDPFIAONB96ncML5QvskIlmPvcfNUh5SbeHZdCj9+FQmsE7jNR1WEeaF8DDs8hgpjY0YIR+Xo1uaw6J1D0vwZ7vbd
Ks1SVkmi22dhm6jIpvSycrc9xeRjGgyTtU17Uy1eerw8Mya2jK61rTEAyhj/jPelIxX6augTh57lShjo8RGPmtRFE4MQid+m+U0Dldr4gYLeXzIvasM1KiAmiQBGwUcq
+gcEKtKDu7GXL4IDhjH1vz+u3fri1Fp6WXf34+so+hJQhBSMMoy23lnOPneeYarUp9DoKoUeQNkaDw3fj9vYtMIEWXcErTmUIOLj5BeiBsLCb4BsiTajugV1Gsoh0CDB
oTdz4tYKjCOu7GR20LBW6MEEkQvp//qXl0h+wvFSP3H3ZfPjRMqhh9oSBwc6k8hJBtDGUw2YjJL+PvW2SYIqcX75aUvr6UpjbuJXfh01SO9dsJ5ZjolSMGIIJCOIgkYI
GcJDVh4Mv6UeL4RK79Ir/6XMNpsqUFhPnoqcQepwCPVAvGdi1sCgUZLMWCg7ySyw/GAicB9buaEyFYGXXrXiXiitbffPq2Q7BpR+gs3a2LbKwyyJxgxiQxGA4P3Cm/Z2
2Yd9nXHs19Q+Uj3uK8qfzkC8Z2LWwKBRksxYKDvJLLCMD5IcrjA1JdxScLlQDJRuV5YYrceM1MM99PTZH3M29frMoqQc9WhEFgO28rmdl66SYt0RQ0Soqs8od1eXCHyM
ZzTYUKnUZeUTPjK2fN/ojYKyv3H1z3wlmAkzvk9K6AM0veT/mjUfRhl3yJqPV+SowPdPCVSv5Oqdd1H9onOzP8XoNfDUXZ7qFesK2KvmNMBYw48volSAEdNJZimY1C8C
20jdaojuFGvUiUp3i/3ZTZdSFBgHVD+wTsoyp152CtcOQR18pLRP29xIJAisYzoxzsHo3iix9PvTfyf+CxEuo1Qt01EVmg+ZCJxPwyBv2Nrrh9LQqxSw6+xeM4CdQKpm
Ks1SVkmi22dhm6jIpvSycnygyASWR6JjKgRDMw5I2hVZLnjEPctdp/t9FR7SVKMNqikDC/IUuitXdYv4rYCCpK4+z38o72UhLHvIZBMav48/aa3juOzDrRHfL3HxpLd2
6hNC3YnDkoPUSlDdqcZRtbbBo4qIwESTVf7i0VMj9egrNyeDrw4WvOch8SPi5c8ZAJp76I783l5m6+HpB3Tm4BVr4+VNVm/oeoB8P76QUnC8+vHJsan27PBsIucLQtsU
Ia8UVg3Xcy0k5hw37nIL8wfScvM3LuYgiVXC+rm2haoYYlzhwKCIAfRPXCJpw4K7uJGrM8DtgVEL4DYPH+coKXOA8i4iw3M7z/SAWTdF1KNrk2UJpa/G7CTg3UUXV1QM
EXfLgORrlF0cfLvRwwV/Gm9kTp9VOLwMmhO4KWv59SfuBnToXMWZzf0Z1ARztrzSmUVOLhlcst/gdAg0Tv90jX4LJoQKsG8m172Dcy49jmlyXvxKu9P2/wWh5ODT4ujM
dj+nRbGNC/v+myjFjx8M8X73P0ew6dA8kUeS/Ihn+z2QrD5iLxuP4/fc8ItMVpp7lNYbRoHcG0eQS5OlBF1VAKs9gdLH0KmPZ+KeRXTFKLkEFJgH5Ks7GqP5nO8FqPxK
Mm7OSOatz925n9mOrfrpCWVkYOlzst56kWNcgI5RxKnCPMrNlhaQVVGvDpx/VtiFc4DyLiLDczvP9IBZN0XUozz2swy4WbfyDQqFrJnC/tDdSUUD9cMhuazkUAWxebGF
deeNY5GKAG1qiqCUCZl96OD+uUHP8iCVihsotUcQdW7GMJ4QHtiIAiq/6ry0Yg9PbHOQn8mSNE64VfX0EMf8JyBEZolRo3pJFuRHbWZoB4yqfb07HARxzCIaGBhsHJb+
Yh8iDKfFqPnolGdYxSzuD9XZ45GN+3WyAzYerR+V+40qgojMdaCgPhjDE5e+HFjjuq/IHhne/emvD9GKJJFaQU94zcV+reDJCankoVbTqCMH0nLzNy7mIIlVwvq5toWq
JBqZI9PuVo7ffYml/tuWF0TgQdsrlPrXmvhgKpDKMCRsyoZ1oMsVikl4fPfhY0mdVLW11n2oeHUu2tD9u3w9djj4ZwvGAk96ckRjzEoUV6Y1gLqX8WBS3xlzRMp3wED2
J1LSnFS9MteuseUGMwUMK45FcjU6w4NCIURIMn9dZL4ETrbFvzyxv4CNCojotCbMwtjwsaEpqZzHCkwW6Ct8PxrGgMht49K/fp4+teMtbedZOPq8JoOY23Chws9of4Wu
8XPIEmlf9LbAv+qpSG4/d2ZPVSaSw0XFyzAP3LlF9xnlL00mqwjItzyHNrEiXN7WfAtnWjgHGPviSHCRPrZTq1fFp7daeIUhRkmfoggacBgaxoDIbePSv36ePrXjLW3n
gHUeoztvbuNGaPj3tIHEwpdSFBgHVD+wTsoyp152Ctc7CGvr/akwtGCBsax4nZa35S9NJqsIyLc8hzaxIlze1p8ctMcbdGSiGSXZngRFSbMuCfT/01I6YMr4rQm+Yyah
yz+W1JkRoY6yudzj4e7jTDv4xCFn2QdRAA+h8yyS7T0GV8lwCa0/ojbjcb8lYJ2H6GaQ3Oa5vzb3oDM0v2yB/9rTMApUhmfq6ZoHS3n0yalTdEGVtOocv43x94WkPs0M
D2by+/IcIJ3jeQ8CrJxwtw71r1zk23wwvxqhMdBce0R74jy6vMFVzcktJUBY0wxkqf2OtUv5zjnWFG55PVbpoBbmTMjGWV/W3Yhh7DcHmo3kNqDYlx6/1qpgFQG13/T0
7jPy+e4y2P0a8Eb8qfEK52ZWLvk55yJIMPuItvbnAF0K8gXpcdMPuNlFTi9Hu5aeNkSVtrEGiLUWXnyReqJvFNpJ3z4kT3B5lCpTEKE2K+veTgAyfuvL/VogC4Z8QuyD
jr1nUSr0UIYkvOglENmrNfb+Ku/6Ca+9aQji5lVowfcjFfpq6BOHnuVKGOjxEY+a1EUTgxCJ36b5TQOV2viBghWhFm/r7eT7vGzUAm71pTrKdkmhOWd/n5cvNZX5BNjt
NXYO+0OBqomkAtR47ao99zSY6+l7YQLgGh0Sri85tyfFVV1GcoewQB1zOBaGFAgoAQUhkXRPMjNM0Db0gJaiZMMr/htYMSS89DyQd17rUqeJi4NLQDf/9P9KyEqgzkDq
Gi0Jl0lYN5pzxQ5tarPbTfd6eCm9NCy8o3zquo1cJpAJX718B/g+h5GQg1/IT9kRzWCcKTHhyAa1wJckP8naQF/VOLrF5rVRKI8/DoH26JmfK0brvszMb6p4D6kcgvPv
PrsOmYDSoKdhbw9T1DtMgxF3y4Dka5RdHHy70cMFfxpvZE6fVTi8DJoTuClr+fUn7gZ06FzFmc39GdQEc7a80hDVBGA+e0AbMcE4nwkgsvOw5RqknQGu+GYGXtwQCX8C
cl78SrvT9v8FoeTg0+LozHY/p0WxjQv7/psoxY8fDPEotusTDUvbrMU3gNk7JH6BkKw+Yi8bj+P33PCLTFaae5TWG0aB3BtHkEuTpQRdVQB+icilHAjNTbYSqiF3Ys4v
BBSYB+SrOxqj+ZzvBaj8SjJuzkjmrc/duZ/Zjq366QkUbxuBUA4MwoZtnJtA62wbwjzKzZYWkFVRrw6cf1bYhXOA8i4iw3M7z/SAWTdF1KOpaDN/EcaRqK5u1MplBCNb
3UlFA/XDIbms5FAFsXmxhXXnjWORigBtaoqglAmZfejg/rlBz/IglYobKLVHEHVuVPz2KA8csvpElqqlHbZOtLfXCIv2ku9q6ca7wAFnxGDC2PCxoSmpnMcKTBboK3w/
wM3F45TRUk8PwSHRp/0K+VXcNuKmhu1fDvRnIj4tHX79Fs2fgAm+LyePPGe5yGTTACmWOIxXuPJHV6DwCt7BJwfvznSrTumMYlS58upXpRDP/UuOtScU8U/eIpl6bOA0
+f639yLGTLignGbH6Ag83+tyhZsQeLaC9Ha2wAxsBQpQFipD5CvpBo/f4i15T/JYfcRCWUTB9vAgQZsnAbf/1k6sLhlGOV5g2ab2zQY3bOPAzcXjlNFSTw/BIdGn/Qr5
VpBLIsZvk2erscexl3hT7QZXyXAJrT+iNuNxvyVgnYfoZpDc5rm/NvegMzS/bIH/2tMwClSGZ+rpmgdLefTJqe3S+jjlRsybgSu+LrS+5K+wnpTl0rWNHrOBMWBrsaav
2JM9/4VlJn6iaX2+IhGi/3Y/p0WxjQv7/psoxY8fDPHivqaTfTV9osqZr4yl3C32ly7nCcOwLL6SjSM0sahdSLz68cmxqfbs8Gwi5wtC2xR3Ky6JhFc6ij6dWPCC2LMx
PDSm7zLNC6sGy4vAxA6EFBzKHBH7wTMnJbBI6akOC5UNPo0GnOtgHTqzw+oaFtxIjuYHq5VC+sfnfrVLbaFfciR2iUnwrGclr8B8RMjzaj9Fn1rKvLMeBkntOlEECH88
1PvX1FFYKjFGI8vkltvBvxkYtfHf8eUd2TPO5B0vGq2Xd9s+SEY7shAN2uhwlyuuDuwfUsk6St3xF2dpcOpZfQoHViSbz40KBU9iyugYGm1LpRJERyOeq7FtI4Q3cdHW
iJ1dYIObEnRCytuUSQmooRWjhKvu8iBLX0Uz1UTLBJbeTgAyfuvL/VogC4Z8QuyDLXsdoRH1eKXB/mv6SKxOjl24s/tScbe3QG2umSXFZPN1541jkYoAbWqKoJQJmX3o
4P65Qc/yIJWKGyi1RxB1bpJEqWxa/LSSaXLRMHj6n4Rsc5CfyZI0TrhV9fQQx/wnoMbVejGJ9RthqSNf/fD7qPFzyBJpX/S2wL/qqUhuP3dXrZM/bNxztd7hKbUvR4v3
E2PIFGobryxuRnmt9ZM+W9eXY8M88bFWZVwfIW1WhOmTkzfVvpim8lUwIi9rGWxz3ICZ2MChjJGBITX5rb6yMALOrQyFtvxzE4istgcE6L5lepALK9TknWi8f7sBGoQQ
LcXQM8mlejmRYKEloOfIxvBOcl1vjBuhLmBSwcp+1987DRnk+lhZFJJO+oDxYUE7KQCjXVaCriffx25TrmlIke16Oeea4iaqpnahKnO0kbZS7IWL0HyAxcwDgcihL29B
20rgLbSpuevkk+04ZX1J+XY/p0WxjQv7/psoxY8fDPF4kUVrvIQEmtGinRjFo9ZgaarpnQctu1R9l3ycie7Q2Bshw6/+azjmMNo20GkkYlkAiFes/0pj579IZ99TPap9
/tUQicsjGvjMSNSkFPZcDpqQwCnz7lNCLi3/fR9/G5QuCfT/01I6YMr4rQm+YyahW94qo9lrB9NuIpQJ3/XI/10OOpKSIlxGlVz7XG8G4COwsUZWjRPYrDTyBaoHkj/o
Tyr5tFXN22uLaImsrvfmtMpRSfdgT3U9g7c1d7SqY+3o2HoRPKNUdVxVqYkyzqvXJfbLlBjB1AUkjiWxo38y+ttK4C20qbnr5JPtOGV9Sfl2P6dFsY0L+/6bKMWPHwzx
uVKt25atEvq4XAjIVo2BKP8D4JqiOULSB4asSs6wDDLCb4BsiTajugV1Gsoh0CDBtD7kSDoc1A2FriV5ZyX9Z8K1xAmSZU+w8pY8FL7jJCtXlhitx4zUwz309Nkfczb1
3EFl5fd006HqbNstQ7vFE91JRQP1wyG5rORQBbF5sYV1541jkYoAbWqKoJQJmX3o4P65Qc/yIJWKGyi1RxB1bmdLNxQXZC4DuYJE92A/Pk1sc5CfyZI0TrhV9fQQx/wn
tE4Ov01J6auoLO1S/BTcMFK36Dy7bTeUZm1eaEPfTAKAO3YZnjpoyC75NRk3Bvqkr0giZnc+pTE2k4lhtKw4+/1cjvxqDH8wkDUuQCKnGi2Kgt1hUiInrLAaTtXVh3yl
3Zg5yV6f0o2kYMP483ZLa2zKhnWgyxWKSXh89+FjSZ1VDOs59IxitXExVs4IDBXlK3FjztIIbNo2sV5vhTAmUsnnwFUeV+nIj0ZSulZAMGf7YX8d61hjiKBASNuth+8G
RvgvXArdBZqoAZKS6dU5fqgCAJMRl9APhz5IbbyEJPURYnR/eDkH881HlmgR8dWkNRdW5IIPQu0sSRs6v41pi8VVXUZyh7BAHXM4FoYUCCgdng+BNvujDCwCyWbz7o1Q
+jGDTlL03/S9WFN1oVCOmPvMaRwfu2CmgiCH1sInQA5RTB4VxnK/j9YeQlUErWD6U/wVoz7Y4QbE4l6IGw7pupZ/SA8VtBy39tymEmy4mwdjZHFlPfycbG7Vz4c7lpwn
EXfLgORrlF0cfLvRwwV/Gm9kTp9VOLwMmhO4KWv59SeR9qrV9RFZtK/zlR3U/7D80OwoCQnTFAtmxZxFl1bWhv/ZcXCYcnOVRX/eZjC15GZygQln0hC9CkJmHY075Dzy
Bt8mf2FYLPqM5hezMZuarpv1gzMJkQ1NO4n+ySJSfYiRuC99fqxREaMHmXgHy8kBysMsicYMYkMRgOD9wpv2dtmHfZ1x7NfUPlI97ivKn84dCfN5kMUIQx4rbFW5bm5S
ln9Xo+sW30+qkYHiTC2CALOYkI2Fy5/i3dTTMpSkKpeAukfdRcMHmpDGiOFUuoLxhqNGQQzqgZFA4xsXg5PcEV24s/tScbe3QG2umSXFZPN1541jkYoAbWqKoJQJmX3o
4P65Qc/yIJWKGyi1RxB1buZLKwWfzMPhtVQEx2xhSvFsc5CfyZI0TrhV9fQQx/wngGJzMjah4qiRum7iolgdskDYhbG89oGk6VnmBkxQBfFH0xmpyWvgYoR8CIZusSF7
tl5WDzzqIQEYMwVoclhC8teXY8M88bFWZVwfIW1WhOnmnibau7bPGdmiNEylqwodwQSRC+n/+peXSH7C8VI/cbKiWFb+4qiHFq7jfMhRK1RlepALK9TknWi8f7sBGoQQ
LcXQM8mlejmRYKEloOfIxvBOcl1vjBuhLmBSwcp+1990Z0Eq85DH516pE1T9+rWR6Nc4DPHFXLd6wqFJmgJOqjMTaZs9+BfVExQOtwEs2ZW7Vdc1bvuHlCG+zsSdsJwk
B6q2M6K9Qw1JF6JHHR0crLlAYjyb9LJXUb3M5DNPmxzKrBlVpYOrIMW+LMmYjXdVbFf9HZFgrBy2SyYz356u8YrF+es5KpgTdsbKostwtddzFihjiJwi2D2tBQ3XD0Nw
lmNiie7sA1LCMt7x53h9PSiRkeMH78gU8ULQQ1GhRon/oppkWiyf1hAds2P6pLSv7bSoZFbWZ8673uTqRSVR1TwzJraMrrWtMQDKGP+M96UjFfpq6BOHnuVKGOjxEY+a
1EUTgxCJ36b5TQOV2viBgnIGPjaum8uYSLNckx1xnw3KdkmhOWd/n5cvNZX5BNjt8n2fT9eWKTEj7ayvSxPD+A8HwhdfpX+cNdFPLgfrfQOSPre5iAX6Y6EKSONF3EPy
lXhsKWIucfck5OTNVIycZ6KqvvO39LqQPdx0SK1+vV/iXTR3LcJTKAS1GK/UrQeyjA+SHK4wNSXcUnC5UAyUbleWGK3HjNTDPfT02R9zNvXWgzRDCgdplboPHgcsj/AF
KkPlVO1UgjZJQZa15WUpkPUgSYHM87G0m/rDL+oRvTAJy39WjlTwqVKIZPAfC6V12KPsAC8XJackk+eY0MyZ9GPVdpY/Yt/bLyeGVNJw0DC/gyFBl7K5f9FFPmiikwBO
D5xzFgNbVlFSEy+XSFGSmXqJb5JhBdeRMzB2JXqJdY0YKvF3LmtUkA2Nylvlh8Ey4jAgtCn+/o6KXpaXTjl1LcIEWXcErTmUIOLj5BeiBsJcKu8K/56ITP6IjhN3MoQf
prW6LyHvTlVnYHEZSx2hFyIWuZNRxiXQx50Lju5h8HwdIYDH6792HVUsHOqymQw1LEz26pTu5b/c0DLxwnvACLbIUnbF5pxzgIrgctsDbumWXR2db6uynUZqF52WgdWH
KXb8ipKjYO/TUqjh0UnBnTjPVMipVwdAUhgVCzlw4rkdTAoNFy3KLsAFKZzjIhoZ6hNC3YnDkoPUSlDdqcZRtdQkuHxq6trsbDWux/7UW3JQhBSMMoy23lnOPneeYarU
qSfx6JBroWpIMDwWGu2IQfFUgrC+69ZeM7kzOig86F6U1htGgdwbR5BLk6UEXVUAC4s2LnxpTs85b0OY2s35eXUnMJR/JX+952TFeWuDIRU5ZrMdl20opbkI8+3fWMMh
7sQpd/odfUrij8rYmrh7tLCxRlaNE9isNPIFqgeSP+hPKvm0Vc3ba4toiayu9+a0/VIsN7woryrYOvMm7yHvKS2HdGC7UPI2AhlyYNzIUL2lNVGQfquBMfxEzy1Al+My
Jr6J0t0X7j4ElFAVQVcWuwXNNv7NcHwx1cNceugkUCPjsZ96sXyZ6HfETN2wj4ZOOl9BPTIGV+S+rq9V5Y1pFNiyuL710KbE7ZI6zgh63b/SCPuOOpV0BrxQirOG3Dj5
NK7LqTlExL8IAAu1IGmrYfyBFd8tfAM/o8HQzj7FYMwx7fM6J/qohsysW+NmXCQqB9Jy8zcu5iCJVcL6ubaFqsTVIItaauHaCTEmWkl1kswh1Dg02Jj24PLFIb1e2N9I
R+sChixFYTT8vEd00f6Huf+immRaLJ/WEB2zY/qktK9SnSXeqacxjIvjjL+9wikR422dTYvnHMIs0Q5bsbymxDWAupfxYFLfGXNEynfAQPYnUtKcVL0y166x5QYzBQwr
csXAGQkJh9NH1f17ibPkijTVnot11dNjlg3Wahae5FepswqW+xJMMCB1nFaU458J8iYFmLbIz9Wh+D4i/j/ZiU5IChHM6KRqspZzb3mIQ3/mjTixyvpwZf+uzWU9ZLV0
oqq+87f0upA93HRIrX69X6mzCpb7EkwwIHWcVpTjnwkH3ivBmDZMU93udqt5MiTVUhP3umRqh0ZHbI5KQaKnm/Qx/dc0Gsmf1U5qYbqUqkC/5zHMt2ywb3/QZpv5rw8X
fboZ6gA2MWywLgQLEIemJ1kueMQ9y12n+30VHtJUow2qKQML8hS6K1d1i/itgIKkrj7PfyjvZSEse8hkExq/j1EizVLA+z1i6BJwRYXUbGzUElEiHRJTFYvB19Lj2mmQ
ACkiINwmRJsxutOVz9rIxMOP2S/y6ltp6gvnJgJsKaoGLNHeQ+SofFKE4H/KDOfpuUBiPJv0sldRvczkM0+bHPHEfVPK/Snn1VfBYcWiE4pGpNVeYVtCqPPpE60QucCc
wyv+G1gxJLz0PJB3XutSp20aoUJ3kK0Sdl4vnmZhQKfDj9kv8upbaeoL5yYCbCmq6CKKo5gUf5t85YUdYBzJ8WCBw9TAe3/kEgAtpkBqqKTxxH1Tyv0p59VXwWHFohOK
vxGa/74GJimSovIQCLTBj8I8ys2WFpBVUa8OnH9W2IUEj+13ZJd6jurxfsLNzVkAd/v9PIhytoo16Me7E9TMImNkcWU9/JxsbtXPhzuWnCewsUZWjRPYrDTyBaoHkj/o
Tyr5tFXN22uLaImsrvfmtMpRSfdgT3U9g7c1d7SqY+0TvDh4XHJ5LWv1oMXgZKWBCGrEZ1Fm2HBdsokVJjjPsChIegnzxbWdxGGHNZwJpgLOrNoj/P9rDfdtASaTxD9Y
f8TCsMZEU0mnozsX248xToltZEj4r3pRM7uX5CLnH7z5/rf3IsZMuKCcZsfoCDzftqtC2GTNu572IIpE76vb3wwmoGR1Ptkm7jKhJYUjD2y4I7W/CGsb85D1Hs8UBUr5
HHmp8/oXHta69rxeIw6fDM4rOLutUhskujKu0P8jKh9Xlhitx4zUwz309Nkfczb1KQDaFBnf75e+Ve/k8g2+/kE2GlQ082vNoSCLUj2rsEOzPxDfumxQdkY//rAxeBcq
a2KoULLq6hypwk0Raj1hjVZ+qLuMZ6QpfDAk2rhlT6zON0Y4YvV9kyDqhGWYhYLMkJ9ZS1RRjHJtNdixg6OtWcOP2S/y6ltp6gvnJgJsKaoGLNHeQ+SofFKE4H/KDOfp
uUBiPJv0sldRvczkM0+bHH6fISNCYDzPDXHS515xqdUaIMR7eGV4MiA+oU/kz/Me92nJRq8M82DXwvS7EUkf83vJyY72yYqWN0pvb3wFcAN1Q5RNf23FdPK5J17CS5mX
NQo89a7qj9/aw8mkKlyIzuQ2oNiXHr/WqmAVAbXf9PShJkde/7YiCScIl/Fels5D5S9NJqsIyLc8hzaxIlze1p8ctMcbdGSiGSXZngRFSbOfGeCvubodaXQC5+46lkUe
PXQGCH03QLrP8JanvasVWQRB6mmdK+wqucK15OuLi/kHpYqGpVLf97j0K2VMEFgmWhEjQH6uHJE/SMpfZtSqmJhpEzIyQnygJD6oU5NU8OXAyOEZfcemQY/ubpKmaogk
OJ64nqjE5ClLY/a/FUKpijMR21OO4F61tttaXZDZb+AMZklYJ7Wuu15DX7OM/XaNRaojWbLQBPPqrOgveHcN6wDyS04lPuVjaEmCXNQu2ZCXUhQYB1Q/sE7KMqdedgrX
KvN2ZH5ZtG5dbgTRGHG4ZugiiqOYFH+bfOWFHWAcyfFggcPUwHt/5BIALaZAaqikpVPdRBoDs6f1jBf+tj8O5ivyGkZ9qFeX9hGM0XzHSHG9J/9vILY/7JxedG1gBtpm
x5L+x0GVRSyjTuQjapVCc3gY2e/zvfZfEWC2A08EminJ58BVHlfpyI9GUrpWQDBn+2F/HetYY4igQEjbrYfvBkPaYZn+AnPy4xrt2vPc8bfEebiArQvLrqbDphk2a1ja
FkBfpRlW8ZHvSZYUKse70RVlb6SF5RvvPuFbVIxqtwCDnEZmo7erPYybD5ft5f/hnXluMaXoiUiYOthwW7QF50M4U52YdYAP3UXaE/tT7VxWUG/uNjRdH7qK/t1f5muO
V8Wnt1p4hSFGSZ+iCBpwGNB/NjtIWO/BB+7EU1cpr+Bx6j8y9DCOMNI06lra77u9eP6sU3JHMCc6Ik+9xTCcE9EDQb9JN95LNxp5/3VhXqd9hBj1rL/BqYm6Ok0pNGKV
vSf/byC2P+ycXnRtYAbaZgjbDh78TL02wt6IeAQaPWoOdBkx9RkWCHPOwf1xMexqLcXQM8mlejmRYKEloOfIxvBOcl1vjBuhLmBSwcp+19/F02ry0CJbaYSlROhgxIBc
xqTGjwpeQVIT5W1YB48txqZ9tSkjP89ao/dPlQqQyleDnEZmo7erPYybD5ft5f/hDuwfUsk6St3xF2dpcOpZfcTKfTDfcjWHRXCzQD0nYNzZh32dcezX1D5SPe4ryp/O
YDsm0NN9chN0mfLOJPfEo/i1V3TXAWGmlB9z5kSBqNOZiOhFYujAbKYR6BT7UWFGSgcR0N5YskXJYtZW/8V3lbniZSs2iCi7ZeesRoIQJFRgOybQ031yE3SZ8s4k98Sj
Fgrgq+jPLXVYWzy5UOzsWbM/EN+6bFB2Rj/+sDF4FyprYqhQsurqHKnCTRFqPWGNoQ7MKuA0QqYWV8/POBUaXdbNmEH9/sPEay4+GRYGXcn4yjoLptDz3kx4+1yTTd63
MAgBDdN9lCxhjyJM2NhIJsjpfSf7SBX2PzMLazHIteeb9YMzCZENTTuJ/skiUn2It7fXA2/56PBfXazYazlogHy4+09Rj8AXNLVmyrL/SGRQKsBccaQX/08Ge35uW2ro
wOXI5ALM7/m2cd7lhtiOc2X4mFqWjKdne5vH6knFPVhiIAye2QBXdfmxAKif+soS2AFNJ+n5vqfUimTumZZlmJOJAOn+ye5V5a/N7NkVbSmWY2KJ7uwDUsIy3vHneH09
vxB+NAXjXJCAGsvFwq3EKr0n/28gtj/snF50bWAG2ma3t9cDb/no8F9drNhrOWiABEHqaZ0r7Cq5wrXk64uL+dlUTsDdbTg6dRwi4HxkQVEpdvyKkqNg79NSqOHRScGd
OM9UyKlXB0BSGBULOXDiuc9QVPztiQs8N/KjkqkgXw3qE0LdicOSg9RKUN2pxlG1lb0MPsnGjj6nIkyO4PBtG52GEeZE762/nZeWb1VctcFYw48volSAEdNJZimY1C8C
K1rIKTB26xsGIxwiQEHduPR2pTEJhsAYQPJoN3+1gXLXl2PDPPGxVmVcHyFtVoTpmer7eZzWG6L00TK3sohLjuQUV0pConEud2Lc2soh0qm4I7W/CGsb85D1Hs8UBUr5
euST3pJKXwcXIxrH8+i9+z6/NV7sZsiV9wAPM6l+7HveTgAyfuvL/VogC4Z8QuyDim8B0MgY5p73sqsXRc/4No0ZeW8IDghfOnsYxfhrp8qO5gerlUL6x+d+tUttoV9y
JHaJSfCsZyWvwHxEyPNqP9lrCiQ50zgFkH4yaE2Ia3SbDp9oJRE/cPf+//QT6CWfnSxuSPvefUolHXbOtrIMIPyu6N8NTGcoy8BoVdqYBEjbSuAttKm56+ST7ThlfUn5
dj+nRbGNC/v+myjFjx8M8VPieNFMeh5JqV/oCO/J7JBGpNVeYVtCqPPpE60QucCc+jGDTlL03/S9WFN1oVCOmNEHqa3pf1PvYuCuRi7wdd7700WrgeHKNlwrC1wC90gY
rVuiznbsfXH4C/plVXABlr0n/28gtj/snF50bWAG2mZlDiGYV/KFLTtX0APgkyBbBEHqaZ0r7Cq5wrXk64uL+QZXyXAJrT+iNuNxvyVgnYfoZpDc5rm/NvegMzS/bIH/
2tMwClSGZ+rpmgdLefTJqR0Fk8rwKvlagtqVZiLopfEYWwCnYZLbY6ezkBdwek/Xjns1mQSnmJNA0IfrJstFFMMiNsGE/p+bVrQdKGgSOaUbPzIDksYhx9Bfj4hB+Wbx
x2MITAJYd/udNEWgpvMKDqKqvvO39LqQPdx0SK1+vV9VPLx5aflbatFll8L++TIrOtPQ+djBj09PnjUwS7YhlN5OADJ+68v9WiALhnxC7IP1uObsTBglVYIjTV8zIOIG
RbjuzlJWyZ4Oh2CS4zsv/6opAwvyFLorV3WL+K2AgqSuPs9/KO9lISx7yGQTGr+PvLf1XxBamXf9B8oLfkf4zk+ghOAKpmGDIMmvi2WIK6GoAgCTEZfQD4c+SG28hCT1
Nw+HQei/un9IfxVu3BFndQiyVRM0wWgd87AEOm9pxJyXd9s+SEY7shAN2uhwlyuuInHQMdG/HyiucfKc3qm4GaWBFdOhminbTgSi053BUEzEcHCey73BufHhbckLS/g9
oinFTQA2l0KsKTzqufEdIxq5vdoe4YbirrR8+oAaPGCZLuVTCm63beNmj+HfExwdRmtEyTQGGu2UqHsgs724Pr/nMcy3bLBvf9Bmm/mvDxefR4YRmfpfe5G5fqPSLicb
mCDfKr3RWWMna83Nb4K9stkx/niARTtdOrk2kuko2nE1gLqX8WBS3xlzRMp3wED2J1LSnFS9MteuseUGMwUMKxOAV9IUpPFTIhm+pK4KJMY01Z6LddXTY5YN1moWnuRX
PVtMfQva6sN/Z4bmHD8u8agaKWqh8NQ55bCgkFZnSq0wg6nEYMgTGq4vSmvGgxFZa02M4Qy6SgMCNp6ySI0nqeQ2oNiXHr/WqmAVAbXf9PRxubeXHna1Ih066rXV7XLs
3atug8HwPFyuCygXoapIjr/YVY+r1BhJFsQdBmOR82MHylW84b7NqGCFOkdEF6TvB6WKhqVS3/e49CtlTBBYJloRI0B+rhyRP0jKX2bUqpiYaRMyMkJ8oCQ+qFOTVPDl
LguX4Er1f7w2rhnJ/22yah+8AuiMFmZsSSLXjMTtRfd+ITxQV1Up7fDiAts6NlhVVQhw4B4tC2RL5cnMoPPoTqt4njYrP/k9+1Kg7D4Wz3TPPrGR47bK9pVeOQru7FI0
Y4Xs8Oh2mcce3aa8nbmaehLeVqsxKG6P0s4QXqefkIkX/Z+flY+YjonEF+PKh0AQ3bXfFUGGfrj3UHU7bfmUvQbQxlMNmIyS/j71tkmCKnF++WlL6+lKY27iV34dNUjv
XbCeWY6JUjBiCCQjiIJGCBnCQ1YeDL+lHi+ESu/SK/8LZLyXy6ICgdhtqJyd09OP0cTvbYvsC4+8v7RtTc/zgwtmOagUSgMZ85ORlKMb+18O7B9SyTpK3fEXZ2lw6ll9
n8cP9erYZMeoqI3+yztsYuQ2oNiXHr/WqmAVAbXf9PTRxO9ti+wLj7y/tG1Nz/ODzsHo3iix9PvTfyf+CxEuo1Qt01EVmg+ZCJxPwyBv2NoRZxaaB3WEjHtZmos2Jwv6
kkmG428ZvAsfKfR7lyvC5qPmBnnuEapmKVYbPtLyN9+ObNPHNWWww9HP87RcNGm4yefAVR5X6ciPRlK6VkAwZ/thfx3rWGOIoEBI262H7warHBs5khHeLLi78HSTqk19
qAIAkxGX0A+HPkhtvIQk9djs0sXdH39JOoIIPQ/uj8qR8ehi5TCI1Oqn2kzmQ6VTWMOPL6JUgBHTSWYpmNQvAgDILO6FEb3ype28bSya8gr3aclGrwzzYNfC9LsRSR/z
0Hu071kDtRdtRfif02TU/f2oOTFLeCwDLhBVbDGxhzglqzziz9nfi/TraK3f0SUfew6VQWLl3tXDlTtCoPa5Lj3LoPcaNskcA4ZjVWZWgIrNiaVOSsvPpDXMjGDO27hg
/+uIJ9qjgOvOM+ia5viXiWNkcWU9/JxsbtXPhzuWnCewsUZWjRPYrDTyBaoHkj/oTyr5tFXN22uLaImsrvfmtMpRSfdgT3U9g7c1d7SqY+2OhtnvKn51WH44Ay+yiuhd
L8gao1S5yGXuaR7pODIBH/+YQg+oOf99dVWE+AuCzKa3f56r2qmScTkqnhWmQIJsE7JJSOu8uCTa4cySetJ8I+zrmp4SXEplMbqTuEJDu1DsATtnWxGOclw2TSb1Fylu
RmtEyTQGGu2UqHsgs724Pr/nMcy3bLBvf9Bmm/mvDxfSKw5uJQC2Vx5iUeAKrysvPDMmtoyuta0xAMoY/4z3pSMV+mroE4ee5UoY6PERj5rURRODEInfpvlNA5Xa+IGC
Xk93YF982bKwrRq9m+PrAcp2SaE5Z3+fly81lfkE2O0dO9Fqk7OpL5oP82RUV4YXIccmvcAwm5GjqdxU/ZfprCLeiD1Iwuyjj2dfzDKZJbFiZtlJ2uYt07kNmg0ExD9+
15djwzzxsVZlXB8hbVaE6QF1yEvlwTJD3pVMsShab1ORj7lYEBfVtAU4J07AEgSWZoXsJ6Wok+hki55v4Y3/5gUnJYalbBsi5Z+ueVT+40aMTczMQWPj1PMT69orIfnQ
JwSLmSvuo6SkOiYgtSlRNZJi3RFDRKiqzyh3V5cIfIxnNNhQqdRl5RM+MrZ83+iNgrK/cfXPfCWYCTO+T0roA+Z+3J19Ly60YYFfV11jEPbWK7+m6Duy800xvXT1WLLx
XssNZRQZqnFMgluTFGUtV1UIcOAeLQtkS+XJzKDz6E5KhrAGA/AfN9NMK7xpmeYeaompCitqZGmighNiT1aHlJTWG0aB3BtHkEuTpQRdVQCkcat4LShfHkUm2W1YbL79
ZCU7D1+Xep7lQ3Gwr/EVfIxNzMxBY+PU8xPr2ish+dDyZwH8x8b3yOR52+T/43VyQTYaVDTza82hIItSPauwQ7M/EN+6bFB2Rj/+sDF4FyprYqhQsurqHKnCTRFqPWGN
p1lnLJnUQS95Zcs9ogNsi6YH7C802CkdXmOyVN7y42Rku6Zdk9kQBDVqchg4/HrKTDMEa4XfenPL1fI3C/dlWsVVXUZyh7BAHXM4FoYUCCjF6j4V5z6HNd4w6t3Fza/x
JZ5Q8SBaBRldM5qo/ddA62OF7PDodpnHHt2mvJ25mnoZ+S4ddfoR0NkWuyDpE40c+ebo1cwagI7TXbjGhngs4TJuzkjmrc/duZ/Zjq366QkODlgN9Tf4uFmVlVOslDOH
0tPSl/9z6EEu4zjHSMsEJ7/YVY+r1BhJFsQdBmOR82P24eR3bS6BSVYXOrIgZa2NBBugXDhTauwwHWQwCgtgJTWAupfxYFLfGXNEynfAQPYnUtKcVL0y166x5QYzBQwr
jkVyNTrDg0IhREgyf11kvnFTiXvUuSX0R9cPQKPXUs/tejnnmuImqqZ2oSpztJG23OzFh4w/YgriNivqXu3atQ5uZzdeb8MOvWheqbgPHBC5QGI8m/SyV1G9zOQzT5sc
N61ZCGPigO4lZ96KDoAmqI0MAwtn27lwZyECBdjWpjMqgojMdaCgPhjDE5e+HFjj2IILN/lrUAlLcfaBZ4hjCtcA1p+2nL+Gk7izcuL3sKcH3ivBmDZMU93udqt5MiTV
TvpWB8lzLpfYfJuxHl8sh9iyuL710KbE7ZI6zgh63b/sQHVZ/8HdCdY3K9+CyeZ43k4AMn7ry/1aIAuGfELsgypBzsWHQLOXV7I6SLSjdNdvmb1dMlj190LA+jBnMUUs
sLFGVo0T2Kw08gWqB5I/6E8q+bRVzdtri2iJrK735rTKUUn3YE91PYO3NXe0qmPt+ubzGE2jbS0J52WKXCAmI4WLHdAXiN0kTWh48Rsu57arIytHlJy+cGHqH09/HcN/
r9yvEq1m66TFwrdEPmrfSFg6YVFy6JYJzJVMoBT3vl6xFl2mQSTsqqQ8XlOOrARsYjLSd9Uwv4ZYKaqsE/q2vfHgSF7od62UUsLd03emcBbKFwS8cpLXnG4Mixt2mg4A
WDphUXLolgnMlUygFPe+XoRBcf+Yj1i2Ef0i4R7g9tyqVXtuh21XxBf9brdaJq+RgONeAw+uPsuWaAMwcuLqgH75aUvr6UpjbuJXfh01SO9dsJ5ZjolSMGIIJCOIgkYI
GcJDVh4Mv6UeL4RK79Ir/wIjQ/ttSw+9m17GSE1cJP57jDABB7AuM3BFhI7mRBhb8BypLVEhKA7rw8PF+lac6lUIcOAeLQtkS+XJzKDz6E4vtmpXAHIx8I2Yy5/hRKFj
WqPHqmnNynMhOK2MbGcNo+Q2oNiXHr/WqmAVAbXf9PR7jDABB7AuM3BFhI7mRBhbmvrJMLpHi3Kgc0WtrPdt7gYiC/V3BP+ZZpwjDsM/MWcvtmpXAHIx8I2Yy5/hRKFj
R3nB9rtjJByMUI3tQh6DRF/VOLrF5rVRKI8/DoH26JkEPyd48Sed190Dw3TLyjScPrsOmYDSoKdhbw9T1DtMgypD5VTtVII2SUGWteVlKZD1IEmBzPOxtJv6wy/qEb0w
Cct/Vo5U8KlSiGTwHwuldfvOD96dLHpffyKCKR0n8ihfmoXP8vtekdmVgNQcE+2IuyYiYfgXgeZ39L1gsjpK6W4jewrV9ljWppTKLPayQinoucgcPjWmqQ6uvsM2KJR6
9XCg0fG0+zp9R6w7hGMSF/n+t/cixky4oJxmx+gIPN9yxCLlA5Ku4dsWdEg/CaiwmpDAKfPuU0IuLf99H38blL/YVY+r1BhJFsQdBmOR82PQqx+M/xi76gIXC0k/Ew/t
2VROwN1tODp1HCLgfGRBUSl2/IqSo2Dv01Ko4dFJwZ04z1TIqVcHQFIYFQs5cOK5pJ7F2bWJyfAioimRsinGPuoTQt2Jw5KD1EpQ3anGUbUrH/Wn87gcVL3QF+d1s5Vt
BwBGWtt0uKWgcfIyWtD2kx/JE8fA3sMWGTNJYa2mHJ1vrK5lug+bwmfizBqIhQNJvPrxybGp9uzwbCLnC0LbFP5tI5KAYB87yHQBtWtTJOMH0nLzNy7mIIlVwvq5toWq
IjAqNKGNUVM6EqLEAgz8piBqG4nqsFn6zKZ0YVcLeydzgPIuIsNzO8/0gFk3RdSj3ygz43c4Q7LWt45RHz/DlBF3y4Dka5RdHHy70cMFfxpvZE6fVTi8DJoTuClr+fUn
7gZ06FzFmc39GdQEc7a80g4Pyg89YsrfioZTmOS51Fv1GIhh+raQISHIRPnMIOwzpK+7F7GTdLo5QynJjkLnVK/crxKtZuukxcK3RD5q30i0ai92wY4UBJ9Z0cznEVCF
wM1WL/DSZWFZwa9Y5Nnm0c4ki7i1C8IT9K/Lal3l2rzHiCT5kL5fy6DRCeeEH+KkueJlKzaIKLtl56xGghAkVF/qKqynaBX6hxdTHDKTYINVn/IXLzSNosomj3Kgjso8
qikDC/IUuitXdYv4rYCCpK4+z38o72UhLHvIZBMav48cS4LisZbR/LUawrKK+sVw+gcEKtKDu7GXL4IDhjH1v/X92dY/YB5oTAgDthjhaBhWomx+R1CcEhB3GT7q8h/i
DuwfUsk6St3xF2dpcOpZfQX1ozfADA6ACNPuUfYbiCOb+H+j047bJFkD7RzpoYCDFwBc1jiAPwvwlVgzXOKWPJVb7pl016GI73qx0LlL6bYqgojMdaCgPhjDE5e+HFjj
eB/L3Y1UDNCLUH9FarShu2n2/S0qtk3yNgk2wZfeGcoqzVJWSaLbZ2GbqMim9LJyEHfM8pPGeKQnHpF732LE3nmP+KvZhO1HHG+uWt8wiC0txdAzyaV6OZFgoSWg58jG
8E5yXW+MG6EuYFLByn7X38XTavLQIltphKVE6GDEgFzkgvnRUcwUkc6ajtAlCqDjoAUcb6k99fYlYievBBeTlW8Y8r/5M8rZOvnN2A6zcxvFVV1GcoewQB1zOBaGFAgo
0YFxXgcWvgUtodwv/97WvpdSFBgHVD+wTsoyp152CtfSTcjPU7SslVcB7HIBzr5W9prxoi7/0fI1RTpWNJdw8TJuzkjmrc/duZ/Zjq366QmFLAjdZsokqQYrwOwFh7Nr
OTravJWzJ37okgPlCeKTipzu7WdAustEWFOyjeQF3ZjjbZ1Ni+ccwizRDluxvKbENYC6l/FgUt8Zc0TKd8BA9idS0pxUvTLXrrHlBjMFDCuA2K3yXB/s73J+M87GaHUK
NNWei3XV02OWDdZqFp7kVy8LQhJt2UajjXAMumRAxw38YCJwH1u5oTIVgZdeteJeIwt46d/+jTlZhwQ8h+3lGkA2sCHjMuKXScYPhTs7grfkNqDYlx6/1qpgFQG13/T0
1ImamesDZ3sG4MslcVUCXDeJ7tY68VogU0yf+TqDw4m/2FWPq9QYSRbEHQZjkfNj4WXLjmU57PmU4jLYA9ZiTQelioalUt/3uPQrZUwQWCZaESNAfq4ckT9Iyl9m1KqY
mGkTMjJCfKAkPqhTk1Tw5ZyMfZsFULuojrXqeaEsumm/1+QSPvHALC5u7jq1aQRosXzW3mUvZgH4+hqkhI8895cwV+SOtqAimSdjJPhpfrP700WrgeHKNlwrC1wC90gY
jbwGnpKWpxgqe1XR7a0sS5GcHkXB9WP4ZuUUAJMIr5yXMFfkjragIpknYyT4aX6z+9NFq4HhyjZcKwtcAvdIGP8D4JqiOULSB4asSs6wDDK6o2gu7RkweDPjbQy/k5xr
lzBX5I62oCKZJ2Mk+Gl+s/vTRauB4co2XCsLXAL3SBitW6LOdux9cfgL+mVVcAGWvSf/byC2P+ycXnRtYAbaZlosW3UCXQQk3RlLOknwdd2MY3f0wG7YGutQ2WVBrKFz
zZ6L7StPDCGyyeO95sH5WX75aUvr6UpjbuJXfh01SO9dsJ5ZjolSMGIIJCOIgkYIoqkY294p1nAAcI+jS+/7bhFYZYqQLXokFbxk1ThZMOu0PdurxsBTMiisvGfj7ZNj
ynZJoTlnf5+XLzWV+QTY7ZfxRy5KlJjQRmZoEnvr4wCwpm/map4hJgso9PFQkFrS4UUVyuL+JnEs++s7mu4IHPFzyBJpX/S2wL/qqUhuP3eX4CUO6DZ09bsjtL9HVIHf
kLO66V6Qrl2jjIXgVFAWy5N15cVzy9kmJOxL2Z64hZocP1SFKnplunV6TbDBVtpFeBMqOxA7A8eE55bNXDFVcjVXrNcXfsZHCWo2GFWT7K2YIN8qvdFZYydrzc1vgr2y
hyEinfqX80qYT6Ien/O6270n/28gtj/snF50bWAG2mZaLFt1Al0EJN0ZSzpJ8HXdx7LjqNwTBQFopPvYPDABctg9VSQbZ4q0BZDGyiojfuwqQ+VU7VSCNklBlrXlZSmQ
9SBJgczzsbSb+sMv6hG9MAnLf1aOVPCpUohk8B8LpXUBiiUh1ouSAxjc6nAogA15FVkPCyV4IvTuwH+m2L6dyrF81t5lL2YB+PoapISPPPeXMFfkjragIpknYyT4aX6z
w4/ZL/LqW2nqC+cmAmwpqgYs0d5D5Kh8UoTgf8oM5+m5QGI8m/SyV1G9zOQzT5sc1bVtfBNG7jjWZb+hnLG52e0gZ6oriMgYoeDuI3soaiwA8ktOJT7lY2hJglzULtmQ
l1IUGAdUP7BOyjKnXnYK14S8MUz6zaXZ0uo3HLH7A1o9dAYIfTdAus/wlqe9qxVZEkDXofvyVl+pnO2dMIsPACWrPOLP2d+L9Otord/RJR8/N9kY1GMtwEy2nxWjK3lr
Dmvb6kqBhhZv7wjgWxagBBogxHt4ZXgyID6hT+TP8x7OKzi7rVIbJLoyrtD/IyofTqwuGUY5XmDZpvbNBjds4zrosYCPy7OI4gJ92HFfY8c+rgpoLojAJ2K7+rpyYcqR
Kv1W04zHway8YetrFXIaH47mB6uVQvrH5361S22hX3IkdolJ8KxnJa/AfETI82o/2WsKJDnTOAWQfjJoTYhrdIJAmiy8Tx2m/yyDOP9doZ7ON0Y4YvV9kyDqhGWYhYLM
kJ9ZS1RRjHJtNdixg6OtWbr1ipBcJe/t1I45HesvMF6WY2KJ7uwDUsIy3vHneH09VqJsfkdQnBIQdxk+6vIf4iJx0DHRvx8ornHynN6puBl9hRCDvhg8T95i00/2AvQb
zcepop3DzzAnYOSe5/niDv4UJ8/+XyCMB6zToyBnORwKJ8X7YN1XedHOgMGZw0THli/FN1TnLwVSCmr2UehsmcOP2S/y6ltp6gvnJgJsKaroIoqjmBR/m3zlhR1gHMnx
YIHD1MB7f+QSAC2mQGqopPmk/n4hEOg3NPzVr078ejzLCANmargG9fF0xuDplR/3Pcug9xo2yRwDhmNVZlaAis2JpU5Ky8+kNcyMYM7buGDOTWKD746CDF0pZI5eiE1e
ElJeb/54RSrFf54PpaOCRtg9VSQbZ4q0BZDGyiojfuxBNhpUNPNrzaEgi1I9q7BDsz8Q37psUHZGP/6wMXgXKmtiqFCy6uocqcJNEWo9YY2/kFMVTZoZUQwnvpZU6TlW
LYd0YLtQ8jYCGXJg3MhQvaU1UZB+q4Ex/ETPLUCX4zKIMS3Zt4JzvHNpgTVqM9Tv/IEV3y18Az+jwdDOPsVgzJBd+dEm1ZjdCxNVPwR0HIx2P6dFsY0L+/6bKMWPHwzx
frDpumURDmCzspS2JKySeHBHJObb26GTSpVN/UkxCR7mjTixyvpwZf+uzWU9ZLV0oqq+87f0upA93HRIrX69X9W1bXwTRu441mW/oZyxudkgK+kgxX88lrVV8a20r+mw
U2vfa8pa5uGqhDVJCdCFsQryBelx0w+42UVOL0e7lp5aLFt1Al0EJN0ZSzpJ8HXdpx1/Q7RFvLM//XsSGGcEp4xsOVEe/EnTOFbs8A9NftRsyoZ1oMsVikl4fPfhY0md
1bVtfBNG7jjWZb+hnLG52SAr6SDFfzyWtVXxrbSv6bCA414DD64+y5ZoAzBy4uqAfvlpS+vpSmNu4ld+HTVI712wnlmOiVIwYggkI4iCRgiiqRjb3inWcABwj6NL7/tu
6KdsndLtbs6RxnoDseGp6AARn1196Jjx7N7ZgQhxiPnqiTYRj3wyDuSl8eiE8dqFXtCvknlYJiMJepXKGx6XPpzwgx2ZwryrteR9G/LXrttA2IWxvPaBpOlZ5gZMUAXx
l+AlDug2dPW7I7S/R1SB37tV1zVu+4eUIb7OxJ2wnCSVeGwpYi5x9yTk5M1UjJxnoqq+87f0upA93HRIrX69X9W1bXwTRu441mW/oZyxudkLP7KMFyW3ync1y1Er4zoe
zXLUvQld8htXCAdY/VoSB70n/28gtj/snF50bWAG2mZaLFt1Al0EJN0ZSzpJ8HXdWOXf0BGkxgqDPsp8l/NLPvQ7E1FOm2u8Vn+rThLF5w3J58BVHlfpyI9GUrpWQDBn
+2F/HetYY4igQEjbrYfvBhOdcpjibIXN0nnMlgWOzLjRcse1nf3xr26+YPtTCqroY9V2lj9i39svJ4ZU0nDQMNsTiz7pXM11GWGkbwek/Qwd2XB7HCDVJUwhl0e3964s
B6q2M6K9Qw1JF6JHHR0crLlAYjyb9LJXUb3M5DNPmxz5pP5+IRDoNzT81a9O/Ho8U/jIOcdiv8fUgv6pqmV998IEWXcErTmUIOLj5BeiBsIKJ8X7YN1XedHOgMGZw0TH
li/FN1TnLwVSCmr2Uehsme0HvEg4pByLxCSIJO6cYo4x4mbTjvVhO/U2umAM7YYtZ3TSnbW8vMM5h2XNJX6BsrISZXwi3UDJlfZyUfORf0S2yFJ2xeacc4CK4HLbA27p
ll0dnW+rsp1GahedloHVhyl2/IqSo2Dv01Ko4dFJwZ04z1TIqVcHQFIYFQs5cOK5XOSGzq9TCgnY4XHS22DhxkHyp0qZphNJEHvscK3QaIWlNVGQfquBMfxEzy1Al+My
jywxHfYksEwxMEEp5fidBPonVugOkGHg474miNlTjNvKLNMVVOQU+In5kCy7wXYHdj+nRbGNC/v+myjFjx8M8aFkxyv4113V5Wc01Vu632XPLA9PGs37fKCdkszq+fpK
lXhsKWIucfck5OTNVIycZ6KqvvO39LqQPdx0SK1+vV+AbcBJMtlnb5glcvKniDwpAOAEr5QiAF18kITbX4/EW3BjAKnXwL2DXZ6Qp9p3GsK54mUrNogou2XnrEaCECRU
oWTHK/jXXdXlZzTVW7rfZc8sD08azft8oJ2SzOr5+kplepALK9TknWi8f7sBGoQQLcXQM8mlejmRYKEloOfIxnMIHfvPfz3WSnROoW63ZbxXJTMMEEUekavlJz3UYHox
G6H+l8nZMSTBmPx6VO2pIT8nsO7+jikHa35Kb5xSwqv5qkOf+tbEMzdDXEwumTaDsSOcMlxeu8FizGDJOyUzCXLd9AR1g1iibIU+yIAKJjl/7R81it03y7IYA+qm6Y7n
VuycfVuK401fX2Fc8AlMuEbxQabvljqq7EF/tKmmCTfDH793mVrRqiBUv0GVPG6XO4Q9pGBWksVFkM6zG5KHTH84nFN9P+h7Nees3SMMzkHcX7Rj8WqGfMlPNk2LvmiD
CwhTJK6j5d5Mj//HI6zEGJg78uv8hjYu5bdSuNNge9PmxVZn9j53VNT1C0Xnuz+pjCjez2fmTti91hyi3PpQvcLzk9wicCLUkQpoPh4dBsYrt7sfFiBqCbeIta2uVeYa
vpO7v06HZhTOLTYCSWKxEzMwBnlq63oGsVEemet0DXkUuHmdI0jGiuOSYIkrJcZNNMt8y59S62NKw3RWWQOLrsVIFBXPmX6qiX/mucnTYBeXX2O1dgAefoAh9Hcg7juV
sFkJOHQIIaF148u9toKltKEPedt+28qvOo3+mn4tDhrx+UuJgELfCDPAus9AvPo58PWGpkXUT03dSX021QUaqiol4JM8UjGjHnotloHG7tOpp8nq1EoVSzQLcuzjCH9z
AJ2DoRlr7inWKfudwHm81VVvAUtMGfMejlTDu49G3ygb6Wof8zIqB1rtP4qzoxQ21TILjySZ75cmUK1BBLgUizuRjQu7AlAEZddoGJhTkCkTrI6u3UFYBygB8F3L5j5b
fA4Hb7y/0FjFk+bOEzbZDvkO4lzkbEqPUgcll/gSbf4t/SOHJXwsQ5Eb6v4SskeQ/TJxgju6zDK25BYEkPrVXotNZgn5TFKd718vUag5bUGwbKPgWMxmOAULCFBrZJZF
LKt+wKuMz71eVbcmW0LsnyWNR7nawVZsyjG+ADQXU00zMAZ5aut6BrFRHpnrdA15f8Ehyr/Jg65L4eaitZ83UADirCr9Z20rJpkPOJhA5v17L0hgLLnh0VXZl1UWbYvD
YuZh7eRVz6oJe/CCt4ZjOzqb6BgGptYH4UilIs/3m63TtBGA7T/sS8p+Koxm3i69KcibyuXEWepmFjED612xWWiwNsL3iHgkb93BI1ddoemmHY7k4kpBP8jRmGoWJd9y
e3sZZydv3v8ljUaV1ylHLOn4IvoCW+T7G89372D2gHtEG8hmKIE3SrEAudFqZ910dVe2A2SQfX8L1NCzxtM8fohGPPPxvGMHK0fOwr5nbVsF6jZjtklT0zKSbRdP3d2j
6b72TCOXBLweH4kiwTBjyHnLS2esGe0+pB0PR3IAcRkdg5sWs3VWEa5vGnpFF61cbYEabBSLTj9ufb9PNHdAJ7C8DTbrPP0qK+m9ciMTn2sn96LEyIVlLWDZTXUFwRKe
tBGepZ84X8sPPjjPtnBI0+aHmoV4CBjDczy4Zrs1juAxd/3p8tdcLxaxu9UoXTsUJr1vqSiOTKxeg8mM4fTc/XRVu1DqJo99cYThzb/wnuh3N7IdfyjbhnGEmL37eRWk
+1VE9GylsYfcBN6m7Qo6yHFLacpgslMw1N8B3ZmdLgRxIoUv2lV46nwjaKpQuR/2HYObFrN1VhGubxp6RRetXMwzI9YDVPnnUvC6OELkilfpEw185axy9KpvIV3ATaWb
Fe+PrHCCqXWmomEVCnKiqluhQHThOC6P42UquuZcdw0mvKmssOx9a+N30g5oyxGoqPcS/IcfjCAtk7IUlGVF+slBDGhLAD9hGAtWyHNsfS6g8ZwHlPwZEWpL7l2ICzdP
2UNc8IoAm0AtmwCqwcMPwj6MFbcSp7LImwxereZw0WoOdyqI4DoqSpLRtWoln+ObcaGmtz6dUR7eKyG1UBUEOCOH57dTB77vwxH+IZRF9QpvVFQM6SWUIJZr8c97U9jR
jWm3/02QuLSOs3+Le73gbzMVwLL/hPWwS3EBDj07zy0qFyA6BlBqSq5yqXx5lsl9j5COTvD7yr3EWWTEHP3dh8qP7EucFWe7imNqju1MJsyeS2hLV5e4eJsStGe2hgNd
z2PDvnJ08sFpSs6ue5EE6YmruBuqSafwPQ2nQ1hvLg7A4t01D0makU/veUvm8OKT79yoW7uiTQqwY3q8V+DGLcoaNrxRh9UDDMvDF/mgivG6qWj4VyoAkWsIcXykZ4NK
ymhJ+AF/+4xno3ex2UmVGbqdy9oLcZml2C+uWN2VkBAj26Ne7LmhwBtlBPuS3+C1ezNGyqq/Mpqjxkuu54E8cl9/mmGYtKedwLtECb5VhE0TCgDeu5z0jXSmCdBsn/qc
rrYIs4cpS7YsiSI+Rrhp89qPgM7lUBXf1GfNyupfK983uS6dvXig4F+pt0/gRZ+q4hm7NohPL6dFYeg+4OKQYEurxVIkQoh2R3bGMy/cexVFeJ+01F8fZF7tMOQccM6G
Q5dj1J5lQ+lpRfFqjauaInJoJizeGncfLaaV8Tix7omoUUj5++ebmKJA0yXySiikMZddGt65TDMejCgAhZB8wqKpk1D0aoQK9nA6Hd3qeQYu1tbea3HvOda0Wz0ra1zG
BrXPxLxDwU3fpGU2ARgCBEbYFO5whEtgUOB+pREMk1NNUNa5wF9JGN0Ttyzoo+MoF1QD9HpJxJveuqNQdUY+xvlKU4WlKheVMeKParh5i7GMZJsZLUH0hxbVmzdALs5c
6370d0y7MLwwgNOiBhK3Yq59NVrvbYP787xD1pXMKGv+XHLfOXo8SkOsD1dlcliocuY5JUyzV3ZEr7CJbcoPPAPDStsbbUVbNW1VF//m4CA9U3HrvkdFBZ3Z2a3juLSG
QLtyiUci6XblVyv1qgxgGMJDhv5a4qiG2Le7vLHvLYTwFY6Q+BAa+1I9IW83G+DlbaiQkGqynVlRBfnubFIZgSHkahPsdOFYe4shTXN7s2YicsLdtCEBzZjXBd511IyJ
VUJ4G6AuGhkCJwW5YzEzwPKSsilq/4RBXC1SXTC91cyrPc7jpAEsiseqOd1SzmqElzBX5I62oCKZJ2Mk+Gl+s7Hb5SvtNKN62dcQsVZNJlvrM1ngsvFzpo4ssyPpPUjG
idxZhdA/LeN3vx9HQUYI7NOrFn5IUwqe0VcIO4ui+5mAWa4hkFliMyJ4F8CsTp11a1soyEqmYF7Htkbu7HD/XFcih5iD4p62FLhDPqVXTVUdcamdtDod1FQf3a6JsbEm
l62ompfquCiD/juKlA+ssgUvKwIU0sxjECax5OFrs6B9lpg5+wAcqVpV8XchrqIPo71jBDYtEfOzPFJebwMANtf2LRe5C9K4cVukfGxdRtm3zI+prf8cbjE4JkVhqFkO
zGDJhtB/CmyvsI9n7NPASUN3z6ICoOmfXaCpZDXtVWsVWLaZG0/rGfTGD/attuVuJ9oqMbPOFwKc5pUkQFvErzqb6BgGptYH4UilIs/3m62x5bASzbPEtegGD+GcA9bW
0nPk2MdexcFEzipL5cakD5cgcVcp37yT/TSjGliBttxG8gLu1AAsB6xQUS1EJZ4wgiX+lFx76BX4GY3S3UTry/HJe4wHaVh1qQgRx/X7/jK3r3pGDIIG4aOourJOGNV4
G1K2bqh/YRu5SV9dEXsJQrlmTRlndOCBm1HTjKD3VIvcoHh+KaNokNp/nXjMdmHY8BWOkPgQGvtSPSFvNxvg5cOkZBzP3f8XEXUb2LOAYlZzbp8ZUKw+onPN96ZGCY3G
AGx+HZN0SRPfotOaFBV6DKbGSwfMF+8uaSusO/YHwoETCgDeu5z0jXSmCdBsn/qc6Nvq75qtYAtshMwfvo1uuRvPR0ZgXu/FmNfk/llb8LEjpHEc3Ca3rbO3hdcDQpUK
AEzm1U4AUe7GUum5ca4yoOffGSaCw1Oq3DpgUTw9Uo9MZy9O0BGAaP5shPILNyLFyqCGN8LK4BM2Tji35mKeg9c8ggqpQj96wM+caUiQckDB2j1lOB9aymrROpnngkK2
ke7uJhUQfyWvRqf7dkoxQ6EPedt+28qvOo3+mn4tDhrK3wpS+1wiOAjlR6E7OR9RcvPYsmbtSJeXNLanPIb+sFnyOVF4lnKtfHj7cV1z3b5eZmiRVQ+nSZRaijFI3NOA
ewWh4vWeoEUo1EcOW7AKc/LWwf27Tvy9eAvqtRcHoSb1bqCxUlbXtdmiwS3PwN6KyLMpREZlW1g3mt7ISOv9/QyhedO8fdO/KfVmyohXGHMqirQ8/pn5yhZc9qEAB18s
sVllQBtRnX6NKDlxVnza23zG8Q2zHGKwgd9eIrYynvjayIPsggtvCQ9iZrt/bkdB3mxgQio5cd9TWnwPb+y8z5YvxTdU5y8FUgpq9lHobJku6vZjvxpZO/UdEPFruFch
S7m9f52vyQyguS01K2yQUpfxRy5KlJjQRmZoEnvr4wAiSmLQJwFxo1YlTWCYB+q0pZfEo4BAMYwINaQjxAixWVuhQHThOC6P42UquuZcdw2X8UcuSpSY0EZmaBJ76+MA
CqFxBv4qDdCt2bvA65SnWi3BVBkNH4vteo4VDkM/R5PzXrG3kJfa2Ad1z7Ei9dD5uHPzQ/5Mr4pHZn2DSkZHqAp+M0Yqg9d7UzCWk7hQOvTsETkAXeIs0syWhaYhEtc4
/2l+sjJVR3dJEaw62Geek5QsOJyLkkHjO4iTxjX+bch0lhZLe+lKHCjJKufHjbI5LtbW3mtx7znWtFs9K2tcxqbJkHGd2MRKixIp5hY7qiV14VS5C/zR9/F5zTQmZxbP
7yo7sR+Dybc2G8tOs1DEjTL+IWfhLGlQZq5V/MU1Hxm9yI+gN1AnyuaKllMxQUu1usr7SNK9VIFU97axevXYODW9qwvHTY8Kjqt1UFmK60U10ZB9yic6oLhABmd+CaV0
PcbJnXNlVNVOwtncw0ewXs3EWKZtTkFxd5wZAQgPX9Yu3oaPoAJL5RYgmeJXNZv5zXH4RVMwu9s9Z+8XLhFHkgow18hOxOt0wDWWWzus76mFWZP0TDRDoOvek/xidXfQ
Ult++v34cSBLN/z9ZP+nq9dCVM8zszNAJW+bOXuMY8pykImh/4G9fsQ/rRXUEiweu2JvsrSco+FUgBKJDUqYPCnQx/+zQaEHJofpPnJvB2V/H7dqWEaB7+MiXcsbldGk
FVi2mRtP6xn0xg/2rbblbr36IiEZ97dy3iFnaYCGE0w6KcV2/8eivz+fGvIJ8J9edLRnOFpzJR6Gx+mI5lB4iNrdH+Lw16zts1hckQrDCrG65Ot5QN9N1asl0iAeLxZJ
qbuwoLcrMEGau20REmQJrnY680pdxraDqruvwcIdr6z3PGDrAA9cZhPqWEy1Vet6H3dnRLxNv+Yr/LgCCuaY9wHkuYZ265xXCb8hjpFQhilF/jwjc1dg2eVA7K6TSdRL
H+/5bpxTLrGo+fuWpBZtedTgSgOqWck6vcxQi2ypOQLUFoNjTbFJzlQX83YVGIm/CZvM8TFuFCkCBNGL9KqPIJ+mF2donAFdvR9IuGrQ2/4Folqy6E5xKoWTYVc5TiTs
U1A/sogFMoemBhPoiFQCDWCzF41XBSfunC5g2naRWm2AOj5ZRu6QuviqVqVhSVksQrPPD97KjWKi36rC7JDmah2DmxazdVYRrm8aekUXrVw1SOhYfWegG+qqqfGuzTj+
7rJ1277mcl27XPNtbYxQx1o/iKDn+8/WrPJV+2i6wyuew4pKpzjMmf0+Xl+eCFuNhCeqTNkOi436d1r16OecnoAZ3TDne0AQjiF/m2V7JBf+xSc+q5fv6rDdW4YpxHBM
2/bKtlshAIdjfLyduhFtRhLIsmBCbehj2KzAx8xfoN7/EpVm2t5pDH+0KaXMLopd2dLKmdm6UbyrseZgiDe+ReE9oz2KzAGk/BdXuDN/tZYy0l2PWZYWgSam3S4VG2Kc
fdpTbNWiLo14S9oWb1oeg5dBXOpySwUGgHgWNtsoy0IYj6m1csjI4HepAZFQhYU2K7LDvbDCgWLJ4dompIXXMMH19HhFZE0T+FXpt7eWcrauZh8XpnVO3HoJc7MsDVSl
DeUpzTtc2fGBrUrn+ThYAz0UwmC4+s5MrxFzY793nc+LtvxIiFP/UmC6kqztTwJ5dJALm99oJlbWIUAK7CpzmLDD0OF9Wjru9mQlfyTfdXsNR3q6sr6LhFOovOlXmi8m
MLAZ4alBq1Ab1G2nLeawGmsvlktGW+fJdVI/DszNGZ3Pdc6y9B05ttk1oGDwFf1A/O56YtBInolywbwnLliEefGI11qYb3So4m7vsVUg7aS1aSzM6Qeo0LYoVazuzxt7
vW8bCb0YY/2VofyvieOuBfKP7t2TDp2ccI/WbkjCVCv/ALDxn0rDA2liWlB5d7+/5j3Ch9ihTR6vodSu3CGdGqpmB/VKu7S+Ay0kh6oSkxsT5JSXuH+Tzg0HXKdEclTT
RaebyLp+wDLB1j8aPf1IUd6RWendouUo4xw/Ztm0qqy8Egs6bvdqpavNrLOdzA2VS6+9Uc/uv06YtmSsfqYtOoFinoc8IraS4ScbVpbKZNgPACD/q/BGJJ8NWWadIVIr
iJ6uXlooteDvwSyxNhc5MKoyamMg8kp3mpUl2OBylf4ah4ByLCyh9rFcdLzj0+PM5fIC4m3ljd5seESbgxudRah8zTyhW1812beyAiyfEzbzWl1OB+fObfFspfx1zcHP
AE4eV8cxnjT3IFpYxkf0tHlmRWph0ycht3Xj0Go2bJLETliD6qiup51y+Jq7AwiTg5KAVWnnaCt3xvxhC/Ws4QcypABRL5m9FkWTg8sx/br/j9uFa9gveJzGbDcc8R81
i+/7Sx1D0hFJIh7QwFSXe+AV133yLX6Xp5aQuxsym2hzL5q6LeBSm0zRjHTQ1ZGrgDo+WUbukLr4qlalYUlZLFI+oi62U4YdtJpc4TA38ZeEB/be7Bpd2LB5SsHNlmIA
4RV5gG0ei3t5gVs7eUGIAXtN6Vtzn/amtfG4HGldfVX8CvFL9nXrqXZvAioIb0/7GoeAciwsofaxXHS849PjzOPBZzECbTJ1+zV2+hrTbs33rUqOOiTSIdhTIMg5HViu
MMOoCZ+MrWTawNwFP1udB1hGZfkgtkztczWJLLqfZ+DDoU3+85vIH9JZl4aJHRqs8pKyKWr/hEFcLVJdML3VzCJ71B7vBICKX69PSS2d5Xv8CvFL9nXrqXZvAioIb0/7
icAjjpXUvWyx6hBXrmFF0I4wUO+TxBggGcuMQEDz7mezd8CVFryZq0uQMMIsi3fiKZvXhwQvgQUfHqeh/n7U4Q09Ep2BtH+5voyv0AgOAXCKX14UP3H7nGDxaOTGPE7U
7lDTnSZZyXP4vvAc0QJILWEjemgTiLDCqFhQjN3tEMdDl2PUnmVD6WlF8WqNq5oiHRQ47C7XClu0JTDRz8SO++5Q050mWclz+L7wHNECSC37j2cKf7XEGO6v/bfa4VSQ
Y/tsX9AGxPYeQUAEaCHkHAQq+zHnHIfv0T6BDIKeLMA1YKYJvbB53GJt7UFWq+O0lzBX5I62oCKZJ2Mk+Gl+s1R4UEvHB5//3ZWWvfY79p5lomjMaQAkugviF9NENjAu
TGHoboghWBH5yc5BnjkVknq8VRUE2hSdi2XygZ4aZEK6FXv96bRm1nHqoPq4EdBE3/xc0Vz1S+Td2QM/g+Oox26NO1hF74o+HsRXZNYTqLNoabdZxsB4jv/YeLSsBeMK
B69CjtjoqJnQ0Ez8mHxb4AqETOKoeMx3+oWz4vXOMfE/UWAf5KdfJ2IzFZYxtHl+eEnlHs9n7QLUH8EJwoc3WJnuGff+yKojGS6FJ5asw7c3Y1SV4oTZFiBY8gAHDcdt
HLeSvmMN3pZFC+4jL0K9uE26Nb/JW9XyIsHnntUSwt8QxPhZTtuh8Xo4VYBUHOX7WdE66Jmcq/BCIKgX8s/IwpmcrdbXJvU9ZsWP9IOfJjX2Beg2n0yImHA/i4I9C+aC
revJdbAa9Pv945vULw6/hsLzk9wicCLUkQpoPh4dBsY8uDUHxxvLyt0KO9AW2lOtRONzhmHjf7WSc9aNrftrjhVYtpkbT+sZ9MYP9q225W5QZ48p9kpXlZesFAo6nTTR
C0EFe3d2r/OcZrVDYDcm3cXCv/ECJHWQ7CVMJQqIZUM2x2wt0GxrzDsJKrwVSfF4ySGIG9IctLOeJlK/3swD7cR1gCZeLkFvB6i1XZYckghXVO/DYPspPJcnrTalw5hW
gkCaLLxPHab/LIM4/12hnl8huk1znM7AfALzoeyB2h7zLJup3x/2Z+xjdyymrXEE1ugwx5FMfFejcTcIEEsgLn/BIcq/yYOuS+HmorWfN1BNkCTtzf5B1xUSdub10H+a
j95ZbKk4SBaXBUh/KbbzTRukODeXPUAEqOxTlLdDJljlHvmPrxVtax8xTsI2QoKJBE62xb88sb+AjQqI6LQmzDzSMCnHzS5bhchJK1BoZ2ZYojP1D2/DHhHjjZNzdsmv
LZOyBJrwC1Ed8VTZgbkS6sw7pZLGWpIqo3shqnjIv8v3rUqOOiTSIdhTIMg5HViuvGbjpB5Mbnu7raI0qwfnKpZvQoINFXxyi0Hyq3999G8GXhs0opJWBxxX5lJl2umJ
6wssSVbxMs4n6fRzCbSpdzVUDA97nreNXPzVV6Oj9/sVxXbHaM/eHh5B/25CWXlH8/fjdSEImMRZPtNGTpMeyUZ279mrbSKYzaSnePRBjunamnQXn6tuc2i8LjNdC4jv
kk2IJfFgJsWi6S7yDB8fUta3707ZG/7sZsHaCyv3WOcju/hLzgxRJs2WGEWLzUCLrV8NP6XakXjvxPYCjOtHbzSo8QKFhSQEdIDfrR3BiMjMrD3VlyF325zE7mZMXEcd
JWWtHh2bWIsuIUvrBAJHxctfKPAMTy5zv8PtpJXwTjtPw+biLiTDcekCNDTCDH7oh1bOt1nt/NloMr/no75IFaEPedt+28qvOo3+mn4tDhp8trMPEc3qyjdk7HjIO9Zv
hJR/jnQ/KGxYMTK9aukOk8svppnyfGxkBeDCFUSANnTpLeuQXAl6wXIXkH4AlBLeWkRXbDXZnhVOEIKzf6B5sgve0YoMCH6zJBUa1zKySYXwPVzNTzgqIiLUdVXETVX6
Txgftoyqk54AMnF1VUjK3WUXp6besMf59yjvZbRw8+jqSovSA2q8sXf7hDY0oJuBlzBX5I62oCKZJ2Mk+Gl+syloJ7iVhOeLA7BMMR3Pm13AoschVtIKxetAdspTsrwu
rCy5YgshowsugfimPNOli7ZeRALREiFYQuWP6oEmBlV8J5xExCMaho9+n5zaRPCCCNsOHvxMvTbC3oh4BBo9augGaC4LbXqFZVthfj6g8HAkWr2yus5JtJnN/0gYm0n0
NzKHqnefPbOvPBJVAGKm6K4XtPOI8jvOIvYueMGPw9Rm/RBN1CSTNMcMV8YpthbMoP4QHzstsmW+gzYzTrZhaZSuo3KQbjk/CtN4N3rTo4+0T040vavi5dWQrSarb8W5
+TalaixlefMOvsR0Cvr8k+aq4blkVorXCyMOx5pSmbvc0fFu8Ro+evH4TQ5IjxW4hxqTw0L0v4pA+5hAU8MTh1IdLtfK5B5IGUCX/0qOKaEUkPz3AWEadI/M32i/Z0wX
H+guzj/uRp8or4p5944GkknWswHg0dptXGS3VR3YMcihlpRQSsJsMfiW0olpskVMFFLuJBv06Evh6WDxgmCT/gUK/al73AF9infHdcX06eTpQhgx0W1HZ8LX4Q4rM/mU
WixbdQJdBCTdGUs6SfB13Qa3k/hi7SD+QvQbn8hoQsxRfAlwrPQrsXmit/Knl+N2lzBX5I62oCKZJ2Mk+Gl+szqdLe9iilj0a+nPGbZCeB+ujsh+v1WIIKRtuUYiYrHs
LM0USD54Ws6DxLEDftrP+xjuBvj8hiHp6yK0xFW3YilPHdUODvnoFGZlbj5Orn/RJ4L7WZ+krIf4sacpz1ScajsVltxv/zJQ/V5SvG4TbLaNlvMc5O9kDDU+Y1rOtHHa
QHKoJ5pYTO69P6PmekkET9pWNARtEkeAin9W6yEcSv6ImEKtDyVPx16x6TshSPDjWB2PZvD3lzcPMn0DLSwyYbQOb6frOv5Pg0U5e+jNcM7YlfYyBm3HwECItguDPBW3
SpclJOKN4kFfcJWZvhgvO6fsbYvX6AGXwWfk3BbwyNrq2e0DH66LByVi3yf1QWtnTRAdM+W8gilIor0S3Jw/I+UHWHgHgC4HvQnAV8SHUzkXkKYMy78L6CaSqcQbs16S
ttMWzRiMyT/7EYt5z3csVkC22dnIYfaxsxqbbPA/exiJzMtSwvuJzLmbXqgbkJtQzQA4E7Y8px5pAYe4KurLTUg3ZTPo/GDb6GC2Tm7XjWwZ0WLSK3A5pVPXi3cyKuHY
iH4WLV5F57C2+TqA7g8UZMpuEKGI7K6VccdPeOm5aYw2HJVosfxx/urXOEz11mWWAhRF9BFInuGYnDImb0+QAMXnLeE0f08/UOPJ1lOnn4Saxf/e8AHk79vvDgIl7r6M
vfoiIRn3t3LeIWdpgIYTTNxOrSEnEA1ZO/JyCxY+CikJG+1oIfOck4/6Df9M7mNfb+5EO0zqmhybyNyClFcyygGX5yhoxWbwqbURz3i/lsYdg5sWs3VWEa5vGnpFF61c
c2qqB3KwskGM9JR06jLzpS/a0zl5eP4tb0stbQfECnspeDTxarUvpytwA4kPahTnRhQdt1aWNCDB9OBygCqiLCxDFHxVUCQO55J9aPMfE2IDfpBAzUwa25BsKWmNewXG
lGdwlSDLqwl8gPwUuzxbVJgZfm1nm/E5xo/emNKhtfx5B9Oqg9icnrVdY125D64yqIF3n/OaBdHmyXaNfeY0gvbNaNWVazyeIAfwr9VgD70LglsHhJ5pEaVOy+X6vrw5
J/h/jACemGIYbNZIrSvj4/QroX09kC64dvfdTE6N57hRNPe0PySvZauf4tgrxjpZAb6XvtVU+WbJ7PIOq9XLGhVDW5oWs9OTY3R9W+thdjZxi9SxPBXgwOvr/FF8FLpg
ORmEajM7lBizG3BCcNw0VL3Ij6A3UCfK5oqWUzFBS7VjXMFtHXSYI5Smu2xCENO/WHnCxa4b+rffHh45yrNdgeYXYraFK7Ix6i88s+bIEHnN9RF7+0DbSJ2FDsYDnf/K
dYykTYmpBGrwAZV144MRJv0WgQ+CE1518HMyRqYvgyu7JMRKsuOOvXXov78Wx3K6Hn04AUTdHhtLtjreAW+kd0isz4ne7Iyn8WMqKS1oEmBVwV5F0+teIPBdkVPUjm7b
HCMPxdmo1PnDyLRwl8E6ZBeqPM3QGDgecL9sPpm/8mMSo+SUIffYsY5ZyOpHCOFZBuUFj7cQo1AsDLWlUIDsk0f9FePaMd5OvUSzUlUoGMWNlyEJV+9S5e3CoNBCmLvZ
HmcEzAtP6wSVwuUCrOrzcCrUTz8BcC6ggiimhNrDpTOL7/tLHUPSEUkiHtDAVJd7dEMkwl90pKI5frK0YpT+Nv4ZJkVkpRTcCUVMvzLdGIeUwy9+Qn6MHg7nl0qTgPR2
Zpkm9AOr4xRg3CI2P6f+kp0bvupPSkv/bkE9dD0OoHLycpnt5dCXP4/9xqLMP6Y5+z7OE6mp+brMxF4notKkBDCxor5E+D63+GjBRpU/r22eU0JJURftAKruacubE2ec
zGDJhtB/CmyvsI9n7NPASR3wIlwk1s6/fFqCRkBchOJsQAead4Yzxm5qoFmscmlxqVzDKnVJwGHoBtki6TY68hDE+FlO26HxejhVgFQc5fupXMMqdUnAYegG2SLpNjry
eEnlHs9n7QLUH8EJwoc3WMkQpPO6i+67PVnNBSaBd1fqvtv1g+f1NlXn0mMtVz5WS/ByNMvCxM8y2NHu9DonmwXIvEK3GCEVDtyGOjpRL/AB5LmGduucVwm/IY6RUIYp
CtrQIXSE/K0RK8Lt2AO0Lo39f0tcShhILrCAvGSUdGXN9RF7+0DbSJ2FDsYDnf/KcvzonnMdUntNnvtldpd+dNmY8J993AVo0sALQqAW4NKIHaxYjU/KjVXfdjOk3dic
ucA9/kYqQ0XugypBlTOZfPRvHHmXsuRvbojCKnYHI3CmFD6iMmOQuQOKp7o1r5qfqPfU6bF+2Fem2GheTCSdULTKkTNoFF8+Qi7bclRAeJhYZWzDbRQ48fStMKsr3Oxo
XjyOVVSZORfh+eEi8rEbAkWz8MiiqbkBAj+YFMK5n8SM/vnUUxKz4ytxi2BZRBSTFIIzoLB8QdsRJunq/r4xejMwBnlq63oGsVEemet0DXlH5xdAeorBnmA9wPAdMBtG
kpL7miVXKn3bmnSDOrKRbiHQRgkOI8LWQ2qAz9i8Ad4VZHowq3ci9hs074QRegFqFZrI8C9NM8Sr/jQ2f9X77MIzwTxgI/sQHSfMsV3/9gnmdzJ02AUbxjhJva12DmYT
kvsUx74E1q6Hw7ql/ZQLJYiE1xy4I8hNv/UgMClI2PEWo1ybQ+PJRK51HSGEhaCjhqI8WQ2OJWXxEheCTpZ9RrQC49654MKR9L7BxQUowOVUdwdefP1WbN67VwJZk85M
kKgtC6obcQUsTL0rf2xK3zGPKIzDOIb+82Js52f2XkSQqC0LqhtxBSxMvSt/bErflh4sUmifzDsxJ38WiLYj15CIBHdWmVdkZTwS8kVtOPkAEpgGLNc/i/imTAj3JgQm
SpuSgb2bxtvqeXzH17p65q2opJFQziQBaqJMdGuEo/HDO6aIO4Teg90pi9cho1RtZaYJJRxPbB9udRjz/6Qwb9ap610vwKh3GMfIKdHQ7EXZvjO374HqUKUKhb2xC5iG
EDrKauVyOeU8+13wOug5vNrPWthYOqx2PjCmoMvxOHiqZgf1Sru0vgMtJIeqEpMb2lY0BG0SR4CKf1brIRxK/uArR7gMatD8jRlRFDgT/5s3nCTBIQtBkfcds9E0DZtd
dbx5ffwoUnGHgzyhOz5KLAc7nt46OfoE9mEU5Jmty5G8KrU5au8kYFEBP5GN92N1Ns+VYRj0vJjm8rcE4ogFB7KsVOp4LrKrmdpDhwdHZIPWSPMNwfGSwaYE742adsv6
N+m0tMknR4/rSzYCKiixNM7SfQtSdKrbHy0vuwmwRW9+cLv2Nb5BG8StQN7DW+p+8N1aPxmevwymdDSlfwHvUDH+wyrq/86faMA1h6Sdt3i5fvdu1tB60UVMr+c7/oRG
xoWCfz6Wju4hCHX2bBVsdrQyAtHKptzG18ou36AocohZE0KbM1YeCNIh60cvuyVguZ8lJB4vxLNfahqIDjsrwX5wu/Y1vkEbxK1A3sNb6n6Fw8ZxJ1R4YP2piSAIVHzQ
6b1Cubb2r8sJ2YgTkmBuLeFSFFcOzUf+ieT6NA96UE8dg5sWs3VWEa5vGnpFF61creFNTydXkSpshgkhurHyM0x042+GA+cD7cY2FxpBEueOUpp4iUm3O0Jh7GLz3Lsz
X+vuzsz7x/kiLg7NbFD5RGWmCSUcT2wfbnUY8/+kMG9Kpprzwbkq2pyYuE23YgF/PtAdzdE8fKferu+GSBvP3kzXbdSsB3AwOuIyXvDNsqG2ZBjOBt87IRYiKFtJpZZu
QgSb1hr5OwlNXbJSZ2/PovHC0BoZwPSRwd+KFioje2G7wq7l3Mwt6NQiFk8v0D3RwY9fcxmx0YyjZa8h36C1kpadMmv/099LaOxoggBn3dVD7DTU4kl8qHU3ktAHrrzY
8K/TzLJFRtCd3LLgEGsfApcgcVcp37yT/TSjGliBttx83EAK8iXNuqAAGPYVUlmMC0snGBODT8F1mLkokoE7cIOU07U6CXAc7xrGGBHkfm1DKhrZhj0HBFJFqPr36W8H
n+iC5PmlT8kx8X18/+XhndaKa+6wcNvIxDjX51kkaJrdlJbGWxWY9PtY/bfc5e2CjodLWT2RNASWo5a5/Dp6/9H29/usgLAxCOrmGwKrch1X//Zge29/WF+BawALPGN0
JryprLDsfWvjd9IOaMsRqM/8aiX/yyM7MiC0ZwpiAcawDXt8mq3Ltq1FCXuDIdVo1u7it6kzhhcE7c1KVrHZLirkR4VLfBnJIeBbViusMhjLUu+e/0EOyYsHY3uvnt11
Tx3VDg756BRmZW4+Tq5/0XgZ2cwBNq32FNZoXiNaJZSxE0LS0FBaw3qvEceD5MnwhUCutTv360gveNXZMENfjvMsm6nfH/Zn7GN3LKatcQTUwCtxyXhdg5Wz6mP/RWbC
lg4RJHJURo8Vq2lktRsF2+tSiGwMYAxZFimjPcxcK3HLiSckDfCWPE012qkER+dtMMgFpc41EsrAVinzgzqgoOKHe+tweeU1TfWcLNuCE2ken4tC3K5MG1Qgr7+RaiG6
2c7g3U3tR5eQvDtKZyAntpAjPnWi7kcKiM9x/iG8MX6yarpCJOpjuD4a2lDfrVHuL7lWk08c+5EJqbLChVZun/pMqexEN1SBkROoQmIN2swyZ9Moo7sLLI00P1fMRkQU
nA5HayiYrOhf8HBTFXq0sGxKVlVH4eDW1Ah1R/vCYO7auVSx2AXXlBHERXk4viMbx9TQJp+uadpAD4xzX1c5KPetSo46JNIh2FMgyDkdWK6yAvZp8Qm3vVA23SNdshuk
ZcFZF4eX9X4du650aJrWvPZUBcKObNSFVYASYbp1U09LxTID79ERPDHfQHOP2GOferaMep6T5+iQeNZY9KMyuzZUM1ZhQMUQuS9t7H2JAhpoyCKRb1mFWWnG6cfL8fHH
hB/GUT/RztaPgTo7bDakbfCaEpwB1mlMLklc5+Rj+iRwPV+qLw5xDLVRL9TNqd1CcG71ll0U1kgxuHqaidtQTnUEi3o5nb81zdoHG0/4nj1aESNAfq4ckT9Iyl9m1KqY
dEzUEaFlSTtLN6oYyMuV1Y1dmbJTdn5xFqDltKKOBK4z8riU2RnqUWADvBmRSZ+qtwthomBXu7uxg1iYAUfgrjMdqnTHEoS5ecYZtvj72r3s/4RYL5DCG5e2mjvQcD4n
byRFvXXqPdLDFQY1ip9MO6oyamMg8kp3mpUl2OBylf7ih3vrcHnlNU31nCzbghNpUB+xXa0fNDZrkwhqVhUkYW2zClvWldWxbE/ZFhDrWrNDdvpnVWONw4Hhrxwr4hgB
o5cIhYEor9JVWY2XLl9i8Gvw4vRfx49Qb2cbRRH+dHbd6zwVTIsW+5c6TDsc5jiCkiRoharyQyIEjmUsRW8fPCeIkE2mkPh5uEyONS6TvkJk8VgW3C3OR9tqzxvyxbGq
7r/MHQzFg7ErUSfLgHrs5iW5kJLoLe4au+DR/gC+pBq1U6cRqKSiSrVvh5piyCZoFsxEQvc52YPI829RsDbftUnhqOBCQJF7i0wSnlTTOUN39jsAFc5TaXjscGVsJ+7j
wktjwfv64Bjiei2QSu1lmp0XISb31Vg/COuVw7gTMKNW8DqghSiPwaRKdGR8cXXFaC9BkR3clGFB2CReER+3FG+zUlARP+TxpK/mFs4UgJuB49mDb5fqR/6JKv8Dn6JI
3NtA8o1iYwQsu1T7+hLacNL+OEZnWjn7/rRl3Z6Z34A9H2mZiOJ+k/h2P2pO/r4PiE3Rp9OVDNjqG0g2MKOphgByYGJ3rUWxSKRWkqkTXBowzTrMCwPa0nUafh2QBLA2
4od763B55TVN9Zws24ITaQccdJm59nu8PoGoPdFzD9mTxXvsG4FoBfB6hEJfp2dtgxdoe9hGp+u9NATBldFd8tTAK3HJeF2DlbPqY/9FZsJpzNgRHSEzDlvlTVx9sQJp
rXpCG9dBpJROFcActtmv8jVJHBXaF0MVsvfT6oXgIsbaiUvQjsukb2BRKMt9Lb8qKKDL9W8h/qWxTQJnRRrV1Y1dmbJTdn5xFqDltKKOBK5w1F4nqng0KB4XWDG296Xw
9hKeVpE4C5xB5sxNGHepe6Aq3ecPQAYO6gIfWyXh1MQjT9bxrprRHz3hS0zA4G9Aj6MZu13/LTqSrvNiOfJe0DDNOswLA9rSdRp+HZAEsDbih3vrcHnlNU31nCzbghNp
SVQdFOsAWnZKwt+0mEG8YwZtYDicfRAna6vHYv4SdBEikCJ4WRGi7cr8h2hm/FlYxHnKyvDFCjfVhicOWDLPn2V0G+F6PbHoa80jXZhTs8aaxf/e8AHk79vvDgIl7r6M
AQBtwd0PdlwNfGunmpih5ViQKNWZQ4m7sAYvrKJdXvcNR3q6sr6LhFOovOlXmi8m3rUyX/hTfUDQ0HR4Oqy1tbJqukIk6mO4PhraUN+tUe565osA8YbVRGwzj4OJ535p
Gf/DFYSUkceNiruL1dNbxxy++RIaBweXlub12Lfb8wzqhIHrcmv01WZfcQF4ZdSc8ivEmHK1wpNnOJ/8xDkrg5PRYYD6AvChH7gap9d6Ud6Q616x6N8Y4Ywl7FX6laS9
Pe2k4mEuvv+IRXARLAUBD0crp2e8NQzoPb1INW+drN9Yd0Son0qrKk/9wat3t3pC8GqN5WTZxnONX1n2QvY/oPtPCtySChEefWrKTU89KBPJKdC/OuPQnWmTNsWeiRfn
y58wzGZmef1er6mjmBElGNgkwfW+J1lI+OHKXxBfogKhcMitXIlWI0ite4zLREJiy1jPIUmezd9DZe8Y5m6aSH7V/5eGQ5MYiXwTMC1EAjHNOCegV75/CIZbmw9Pjv8X
/4xnLOdEVW6N5GNCIzfIZewd4DYsJmDyDNvv8Kzz4wMknQCvsjoDP14P5H/HLk/TwqgKhKx1HIcULS4g3iB36iPGwV0gAHfAsBQRSqYRg9Ug4k2dmlM8wsjj6qCfyR04
adeVrGEPkkQ0m6+9sPfI2WATeQ3VbA36ttZE1KKN/d0gt8h5NAzHqFhIY++DKJ+q8GqN5WTZxnONX1n2QvY/oPtPCtySChEefWrKTU89KBPJKdC/OuPQnWmTNsWeiRfn
4BXXffItfpenlpC7GzKbaEPbqN0QDnow+8j5BayNcGUt0BBSr6EhAjFhINalyUTHVvA6oIUoj8GkSnRkfHF1xfi9S1fVG15gl4bsb8w4ZKw4S9dnU7k9XwWZnsKggH7l
iXnIpl5rV3A7BWz2tQURyAZHiyux7MajDZYCjyG6oFQnF+EqPxVkSFWQVVvs5Zv06PIlKHdr7MTk25PtN9BYbUPbqN0QDnow+8j5BayNcGUt0BBSr6EhAjFhINalyUTH
VvA6oIUoj8GkSnRkfHF1xXjyN4xV/qG0jvGFgNUFqQcf6Zjjha1trKH1kMJkc3pLdCwvTg1rR1AGPaEoPMwl7Ou2VDSGuWSGuO6XTN2wlneojHI0/NRw/gynT/ogaYnQ
xxhs77dzx4VomxIg+jIXNh5kgQczDlhYZoIIsxo8tHuT24eZynV9ASdtKPZoaZxxb2FbiBQeJvBGA/31ryOKPi/CKokzbO7+yO4FKrgF3dOojHI0/NRw/gynT/ogaYnQ
xxhs77dzx4VomxIg+jIXNh5kgQczDlhYZoIIsxo8tHtD26jdEA56MPvI+QWsjXBlLdAQUq+hIQIxYSDWpclEx1bwOqCFKI/BpEp0ZHxxdcV2BlMEwJcRKNSpMTVhy9zp
Yn1vS0s/SMYcbCx5Qe1lE1/QkDXKlbhEoIit1MJivrprJeOUN3vY7L5+j9YZgF3CKY78bw42xEgBB9djeJuwtvt9hDRe4hgfNY3kbx+p0SELhwO+9VOYVv/KwS7kN2yH
5j3Ch9ihTR6vodSu3CGdGqpmB/VKu7S+Ay0kh6oSkxtTlvjwy0XJ6wDWLE/CzpM6Hz4JQB3AqneLRRmUoeflBcXoCp/2BvJaELvya2FWI7q8gFUc4GxIZwf/TwMAniCH
SuwnfrFbhGdELP53NAGpk7DIq8ef8jn4tbgUSvkcoxnwao3lZNnGc41fWfZC9j+gyYUUHxAUvT6Wrn+d6phLt9GPbVjows9b2zrp4Jp3V8imh4aATdNZKofNFJpSQZKR
iXnIpl5rV3A7BWz2tQURyPz0Rj8YYZa/R2Ir2m2LVKZGdu/Zq20imM2kp3j0QY7p7B3gNiwmYPIM2+/wrPPjA0lUHRTrAFp2SsLftJhBvGMy8i+Uo1N9hgwDrR0VUglw
vCq1OWrvJGBRAT+RjfdjdTbPlWEY9LyY5vK3BOKIBQen7mPN3n3vbxrh9R6TyuUQTDKAuGKozhaFzNp/RWXDWb7mXeXIU2izFzbjDPEVLFLTc9heN5EMfZagablW/bjj
mJoP9e5AOySIJfHBOokwwK/ULOZH2TQeVwlQ/mSXLhmlRQb+nrvHwqNIAKiC/vrurV8NP6XakXjvxPYCjOtHb8pSNHxGLAyUXOxZTmyJguSW+ccF8F+I/ICJ8UX8WV2B
XwvencjsooUsKMw5KyjM7zCOURz5oFxrW+vbaUuRZiIy8i+Uo1N9hgwDrR0VUglw0fb3+6yAsDEI6uYbAqtyHUKdBB4fRGuzMywJ/E6DXikI+KIcviFWLDV05Cv/JIRG
I2RFY4AWfU1pjx+ctw7c9EPsNNTiSXyodTeS0AeuvNh+hIL1qDRYeShnUzo//5pUx06vjolDZIBIjfaXw3kzP/EpESaxdFVXVvGindNMl6xmGrfMmfemwDE4q5QHCxSq
9DOYclc3Kgg6ZmLRdZzVlEIEm9Ya+TsJTV2yUmdvz6J+hIL1qDRYeShnUzo//5pUx06vjolDZIBIjfaXw3kzP8KoCoSsdRyHFC0uIN4gd+o6o5J00VkHarlQTUJFvW7N
LSw6Ejt0sH2iVNJmu7WzG8g20IZVbK+BlhmCvm2P2Yu5ApvLQbzkHGvSzDBzoa/JBxx0mbn2e7w+gag90XMP2cUp1psPEqn3aI0mD8xsj/iTb1kjBRNM+GVRtL8e8l5t
KxfM1+R8NCRCQorBqC/ApqEcIaUxSJO82/599WfhHDzzLJup3x/2Z+xjdyymrXEEeT2/yUl6OFdMQ8D3TJxLIcaJap6+1Ea+u1153oScsX7xKREmsXRVV1bxop3TTJes
JB81IRzQzA9uWjBLT70IZAuaNQGLch3Rou9WDuevCMZzSnxy3f/LepceMP6gqU3VUdP0vwS8crsz4FGGRZHt15shXkZIjMpRFhZc8fnNwJtFRWnh1wD9jR92gNnkOnr2
yNQeEZeF3npSPt0BwUeMZbqOhMlyDX48YuWgGYXDoHfrtlQ0hrlkhrjul0zdsJZ3wuk8G7fdJpyy/c3Jd0jVzhQoit2WAOkxKQbV6cjZtDkeZIEHMw5YWGaCCLMaPLR7
Q9uo3RAOejD7yPkFrI1wZZqTuFs6pQv1qt4Ia/c4wkVhKRmh/hBb114zswOPouJ2JJ0Ar7I6Az9eD+R/xy5P058Fmv8wB0QHJA5JC5Bvt6o2qlKPy573AFOdevYEmeY+
lBuFlqflEJo4JCyA035507uoy3Agbyd1baqTjWRGn49qbORd6+P3jieSGD3QPgx/wKpiHZSst52frckMC/Z5yBn/wxWElJHHjYq7i9XTW8dvAhFoT019G9rfeto6wZ4I
cLV3vWubh6rtdWi6+DBlrvi9S1fVG15gl4bsb8w4ZKwGEqxYw4zEwW6pr40hAE5btlzbfD8I/nGSO2C4xX+eTou2rH2A1Akkh4+3MPc+FPJw1F4nqng0KB4XWDG296Xw
zSjLr0A6bPBXaCzpWMVo2mW6NUeREGea+pwFW7ppor/T2FjdKJoj0JQJsgyVVWE0I6YAY1pXo56kuxrgO2WX3Iu2rH2A1Akkh4+3MPc+FPJw1F4nqng0KB4XWDG296Xw
NBR91Iyt4/ZNx2rm/dZdLRPeXdoCUtYeXBrEFkT/hdMtLDoSO3SwfaJU0ma7tbMbyDbQhlVsr4GWGYK+bY/Zi+6/zB0MxYOxK1Eny4B67ObOKECZCrHKL3JJYP2es3td
fnC79jW+QRvErUDew1vqfvDdWj8Znr8MpnQ0pX8B71CBIDmjzq5BOyntbEirb/+lWHnCxa4b+rffHh45yrNdgbI4Af2a7nOHbsfdWtkSx+UQ3XTjgx4FA4MPDWjxeeNC
CFlsB45hkDvLY6Xc5vA/4MEGD+8MgNirjfUDN63W1+S3oJu5qEyjtmIhgxknahxM40uLAIymdEhl0kZ3CQXyIomdtZ4S5p3pCxmwvJrorS8AcmBid61FsUikVpKpE1wa
MM06zAsD2tJ1Gn4dkASwNu6/zB0MxYOxK1Eny4B67OZ65osA8YbVRGwzj4OJ535p3w3FMtqRkyp/rpWnYPi/vtaKa+6wcNvIxDjX51kkaJrYF1wDXurWj73M8U9dLOOl
u6jLcCBvJ3VtqpONZEafj2ps5F3r4/eOJ5IYPdA+DH8ost/Z4WkcaZbwsBRivMyGbbMKW9aV1bFsT9kWEOtas7lBywzu7teTdPT51y5I/rtm96E8/OO/ECafThQnVV/8
4IuYMcUjyvv/bX022gGYLJJBxr86hln+544t4Wf9BfA9dzDSAUv7HQjxAA3Y4isPwO56cYyJLrsoMIrdvItaxprej5wXvOv+KppAMCzPozURXFmzABMgfK9QwsgUgQwN
lfg56btW7sWJPST2QwsW4MmFFB8QFL0+lq5/neqYS7fRj21Y6MLPW9s66eCad1fIpoeGgE3TWSqHzRSaUkGSkfqkFprF6HMh1TB+K8+UyJKfm9dkCOsoACYzE494YUMK
FCiK3ZYA6TEpBtXpyNm0OR5kgQczDlhYZoIIsxo8tHttduVITJruv3aqc5RujLMzL5i8HY3Ix3Ok64SBGtVmjR23QSLE+/ewUqbyol4fTfi6FXv96bRm1nHqoPq4EdBE
qipd3e3gKit785SVKmrYpD6V3CmkLVcr3z/yG0tFYKtOchzQ4JNfop2sd3MbTr0G2LYzQ2im2O99oMk90l84ESa2kXCOjHx4j0BlDtPkmZT+CJgFiFUVl09nsVzdNFc7
2fCSZiP7TW0qUg6+6JtnnAK2//I3ZQlw25iEABuZASA96sNQEddbdKGX73b7Wb/ZqAiFsBwMgBtoaRm3YtERU/IfPaRLobsugcUouMc3ITUNBDbVCjsjLY8o/+oikEZo
HzgDPPBhlpWbMjaovAJMI6jalQ0J8JZrP2hgYEQgG/1hVCIGsu1q5/5GJVTV+KmejkcHp9eZeO4AX6cVTdC7iASViXzjJpVN8PvaYD0ZU5XWCeVD2+Qqw0EWw/lbekU8
ayQ1EUzHkBaF2f03nHHcTEwuT3bjR8OhvnBfOnNyqaDZPX201Lgj+MppT7/tvaic8WGpcAZ1HammM1MB9eeNcwnU6a6o2Ij2Gc3vU7Ey4A7XlrNko5wFYpqrs4SxCFhL
VLtOBSFPTuSVSuWE53RV4vREGERsuC+0b+TEbW7Jlf28LFUbrDvUnI8UKJkk5GXed9nNN91hhVlIWjy/zEHOSy9NPlaBdNKdZuED7eHGj8bFLGtej9wPqqQjZEzn93T4
WqgE8OKwsnab2vLxVvgFHaaHhoBN01kqh80UmlJBkpEQ6+xTpVy46S9jZobNrIJJZuwx39vDciPIv2+YssY9Hg8kkMCSKfxnVrmHasGTcoVtswpb1pXVsWxP2RYQ61qz
o3U25NEIjmSLrPprbYrq7P6IduTH3SHC5DdNqMjhmfZk0snPERZDFIWokRwJxZa2mmUbGc5nE8KQqwWZ3drXHUVFaeHXAP2NH3aA2eQ6evb3wjjGAZjRW1z+EDjsT7eU
AQSfPquL4q7AjObfAaJ5geEVeYBtHot7eYFbO3lBiAFnHXt0195sgpI/TPelBiBIVCcbLCEly16nmdXM99IM5mYso6LQZuUAjtSRjXBHYMF310Ecyq+YeHb8SZa3FLc0
GJwoI48tRv6rCgd4L5wP/TZI820OJ97jSgpsPOdBTY9WG7mfgYGWd3nuKw1OUxy3M7k6taiO9Y1Ym3sjmXg9uPpMqexEN1SBkROoQmIN2swEjMafaS2RGS/DsciMpC7M
zCrOmMP9PtPMSsvDb4hj/pZApYm9japD+Tww5Bbu9wdQ/TpTK51+uf50qP0Ey66o9hKeVpE4C5xB5sxNGHepe0g3ZTPo/GDb6GC2Tm7XjWw3vdJCNNf2eIr6Je+nHAfP
v0KtF8vPI5m0cFzKwpbPGP+GkIKGG+35IeF5p9TjU0En2nGCS136AQq5XtCZ29PBB+20mWam6/AvOOfN/mwu0cGthUqA2akUbNYwJyV96/hNqy+BU5tQ3qoeGCsGFJ0j
QSyG2rbrcT9FYFi4DToDzNpxWec5AvWeZxkeOrdaMP5Nzp0r0QmPM36MtmJXa6P2+TxSxhbkps3ar8f2leecWDtYFZgqybwT1TCs/SPyZIAHCYNFUtgIX5sww+lelzbY
qCoj0vOAadFV20GxzrLo55GJbv4SjrBPWtjlq+SzwuInDWpfSAHoyIV+uFGcElL+3w3FMtqRkyp/rpWnYPi/vkYwcjxoOoEKjSOaZHXi7nV9NrVkvm3CDgkRuts58WjY
xYcd/nDS0pwWWsOg7ItznZhy9p1Vv7b8HCK4cxENliu6cmRXz0jRjUDZJpeWriVbiTQUSRNmuK9lP/oBJ1Js3UPsNNTiSXyodTeS0AeuvNhGDySmfj8konTujqUk5wyb
FGOCPB1uWkOOUawK7NdG+5vpma/4o4SdN+VGP8ou5b5JWEy3fyNfGDx/i6h8b5RfjWo0w0BbcmhP/fgkT6f+ITvaLvVdDBNKCvWBp1sz3tbKQeXtN0124KMxcfa42HP9
zmhHYjYrWLLO5EHpZPREXtSGfd2uPOCf37sCEKNkQUt2/yst/ddPQpeaDI8CZ8n0IgJgGux37r4sPfs2+xtb4jhL12dTuT1fBZmewqCAfuUQ6+xTpVy46S9jZobNrIJJ
wQYn8YrTyJ9ITWW4n4TSMhn9/oNNHkEHgu51bo+vctEZ/8MVhJSRx42Ku4vV01vHUT2MfFYder+d1Q9mU6tYIqaGlhsErD1ydQUh1bs5a8KqATxbL9xvekHFrJ3wbJss
FOkHs3pCIt+PSCgQxf6CT/YSnlaROAucQebMTRh3qXtIN2Uz6Pxg2+hgtk5u141s7nqzAxmPD/CbY0W8cOik0Bk736bAIcsKh5bDj8hgL3V1evGnbgUDMglbaPbgB6oU
fWc/3c9KOH1VXj5pUKbFscvsFOUFzdHAiL/jFjmHJNH0IY8driZh3YMkVsLTwyxszkUI5FaC9T7DdqvglrFq4f2CXdBYSdcXqLfdXFQ/sbJaqJu+j09sqpDnl3gSnXr1
DUd6urK+i4RTqLzpV5ovJpYimYOWQGdlME2CHQZNK8omH9jz9K+2m8/HPOmM/gmJfudtR1H4Tkb4/4FA4aWECImMAIf28FT+XkvTfcS35gxVm9QFYz0hJLvSVPqBA5zE
NuwAHAYnRP4PPMijvmPdkAvS5ZNbWLi2c7kHwKs9c3hfDZwBaRuSi9SnnDmfmkZ6miI9362LMLPNZZ9m2lLDRggczAA3jHlp+Ca9jwhXAyKbs5SnKqv2qN9897bs7HoC
961Kjjok0iHYUyDIOR1YroB+FdXHXguSfloBVFSZPIqVpVKx3ImLXpZdwpls2CJ3r6BwoqQxDzXh2nNUGw3TxSwj88ZYYbDcelunFulr/fDvEHzRvTMkWyQb6UEwtIAK
j5MIMzRqIaWPtTY/5+5Ixc9CTMpav+Up0bsi5JRs5ko712WCVXDEUzcr3vJN/M3remDvDVhwXqe9s8tdY28RbhHz1QzRutYFaFOwPlR4HrKqZgf1Sru0vgMtJIeqEpMb
0uwar8UbzPPHVEUG8CvD6TyVRJb8rQhHnUDY66HcmlXoFv2sAxqXNNabzLd3Kxx0NgNkO2j4hwn+GCsY1AOMUR4MbZwJ0/rB2DfaDdvZq9mcXq5v8qxtN7qGePhorqIm
jWo0w0BbcmhP/fgkT6f+IaSzvx3Xs+kZgDRboYPJD8Cw27DseU4sD37CTI6D63v5HL75EhoHB5eW5vXYt9vzDPnXk+jvD7Wg5x2LV3fQP+MQiD/cE+zKudeu86wp2/Cd
VJqDarvZmR20nPQRERYhi+0xGldS0WUZCxLGzFUKPRPp7NQLfygvc/bDDgUeGOMGCVLdMTzexQrD7q2wlL2uy45N5uNsWOY9e3k/vhdOwGDCJ1Q+EiRcqN6nqCIXg38t
9YO/2viV+HV1TZPU2Opt++a7AfNLYKwW5dVBrvY2aXXedbJOTZb4D2XKIPvx84tLi7asfYDUCSSHj7cw9z4U8jOoitQKT6BZgM2FZKZn+zUoUcO/GVp2UFXJ+3r8zHni
duoS0dU+sY1WxAnsh1vwZft9hDRe4hgfNY3kbx+p0SF7KN99izGjLzq0YLYuwYXfAQBtwd0PdlwNfGunmpih5foVZ2UePt7YU0rCNDLxYLOavjO0egC43Q2npyeqsieH
1opr7rBw28jEONfnWSRomq4zZzIprACQgJglKG0nQ1V1y3LUv4K4jWFn12STbYqitmQYzgbfOyEWIihbSaWWbvXhEmvuMwdxevBFc/aTuAoZOr0GpwSqtIKrB4QwcYzt
rwrIZfK5i0ahI7601DOZ6whZbAeOYZA7y2Ol3ObwP+BrmAfboBXyeljr2QiWl2E3C0snGBODT8F1mLkokoE7cIOU07U6CXAc7xrGGBHkfm1VzZoaD+a4UbZFETCEpIrw
H2w43Jlj5ghjaalZUplaYSP05a56MvIBSmnYI91duzzlVbd2otOjJPgXCAyIHSwPbdJQyaRa74tZZEbs6pyDnVjGB+JslaEr7GwHdJQVc7O7wq7l3Mwt6NQiFk8v0D3R
ROjw3pU61h0CJjZloz0gOqoBPFsv3G96QcWsnfBsmyxLOb0LYSR1xqgaBZK/hi7OHZ8SO7VbPkYgAOX6pElMK5i+BuJQOtotBm1LNVQnikNUApft5sRNf+5Aghxg8jdJ
IEE1T9QwL3P/oUK/VnERBPdNOj0Kk4dZU7DKnJjgXa9shs69UmKzkpJs2nuR3OoDouBJ6l6/QN/2/OsgUg7/M4BSUocUX7GEqbRWUlQVi+lke3Qms/e1ynmeuFjk3n6N
vuc0o8wIY0gVIGBMpAf9O5PPvlBQEqq3K8Q1M29SjbgcPUIpv9hBh6iseSgD8psIC7gyyL2M43HR8ff9ltDfBkvXHaUbgEfhjTVE1So7kBow1uJoUrBOWP/DHLjhYDb2
MM06zAsD2tJ1Gn4dkASwNia8qayw7H1r43fSDmjLEaiFX75ZcqJAjZmQI52URHuVWZmP66vaKfxsrzuA9Ch3dnEXtolXaSv1alM1QWgFaairL2dhm7L7tFnW0O6WVBzF
67ZUNIa5ZIa47pdM3bCWd2DnY8gzlAvqocPkr5zHtB/0gfRkCmh1JR7vf1Q3I3/D9Lih9P+smZ2TxxsWRL8fqUVFaeHXAP2NH3aA2eQ6evYmvKmssOx9a+N30g5oyxGo
69Sn1f935RmY9fXXN2zpISe7xkFivcbDCIkOWzxtlY7zbDgRpfsN9D2w58ad4/uKDAQNSG4z8Jq7+asdTahMvkLD+2SqEdf0QTJpd0gpcGin7G2L1+gBl8Fn5NwW8Mja
JryprLDsfWvjd9IOaMsRqIVfvllyokCNmZAjnZREe5U6D59HCFFzvQsmD4Xyu18lxhuGt2Kgp8516mtQ7aMFVUZsmnhtLctfTgCR53SMu/L5uIa89ITr6JGPeVedxgYM
DEj6c9gJ2uqmKuCghrsKq4HFQg8ykhpjw4/m4lFunKcAwfjxPKoXGUBAk0tETAHG+biGvPSE6+iRj3lXncYGDJPV2p8qySF/tWf5hgjcOXv2QSEHjCgJ/7xKYYBTP1Zs
psHHwXrBwij9vf5k2lduOhljaHfncGTdh1PTOGVaSGEsej8XZLelYtIkkyOOTo8FBubpSVSy3vWxe4LrmnIlgia8qayw7H1r43fSDmjLEajEjLqIZRPwfkkCt7tHbl3e
pUaowcw1+8I+XTilzaO0Q7lJn++I2nr34CUDxN/37bvXfwmavFUpEoZQfYCyzAS6Zx17dNfebIKSP0z3pQYgSJ061PMHFXTtNO61JJouO4pXfU3DausIxILYlQpuW5ss
7QJULJrXd4uN4HIolWcmvEBEAsJEh+NWJGl4BZnddS2mwcfBesHCKP29/mTaV246H41MNP+KklrNKUbhiu1rllQbATrOe7SEzaiodE1uuIPTma0401444/gjwFPXDxbs
MSWdqFEk4PLJ8mcotMwlulr9r1HlGwveGRdOy9l1fkAfjUw0/4qSWs0pRuGK7WuWIRk4R9fLj8Cn/XT2WVwrYZZ3iowTGXVvbdTg2NUYy8tj5WUF6XuVbh6ykUS5Z9Ec
bAvy/3N4bdLHXTtDdstDEWcde3TX3myCkj9M96UGIEidOtTzBxV07TTutSSaLjuK82w4EaX7DfQ9sOfGneP7itfrXR9SNqaFDoSCujoqd/iNwJwrrVdEN+a/RDebdd00
Zx17dNfebIKSP0z3pQYgSMv2ECcLyIMYOI6N7f/AvW16nG5LMPj1gh3aT6xeNMpdlkClib2NqkP5PDDkFu73B54J1uaH4+0eZ25oZuVu8Iv7C+auepIViAXUJPXKNSZK
MM06zAsD2tJ1Gn4dkASwNia8qayw7H1r43fSDmjLEajZkwrnvgYMcwxcjCdytZuwuKq0GQ3MFrow3LsEfhVKFSa8qayw7H1r43fSDmjLEaiwYmMD7c2ZrfdufBestamk
QgSb1hr5OwlNXbJSZ2/PombsMd/bw3IjyL9vmLLGPR7yVYUHw7lccA9EweHmI2TE61f3EbK0KIF0xNeK7LVkcOHPD0+aa2R/Qfo5uQJEmW9V/KGbwULBrwv4QOy5wrpr
fFCROi8pQc+AkgMzLZILa4oRxWX2jUbDXX0EW6Z0FC51siXEpye7BR39rSreNMDVcMJlXycnvpHMbHg/uMIK4cUp1psPEqn3aI0mD8xsj/g/PqQ/713h5kkn5IixnOpP
4tfYfaZei1zguvys+5NVB6Z9xBcUjcUkJa7THvE7EcCDliNpzhSg9+stpi3f0pMLkyPogYo+nkr47hywQ660do5F7/StYekJXc7qw5wp/KIA7uucX+JRAG+lVQXZYRn0
okQ9X7QS+sZ6ibZJRlxVbfm4hrz0hOvokY95V53GBgz1GABIjucUODFtzDDD5bIIAe3HDDreuem4YWxbxCRCNuLX2H2mXotc4Lr8rPuTVQclisNZBNwo9BqBzkUiyTwC
mB4vtsJvAJtIfWGhkLFzkgfttJlmpuvwLzjnzf5sLtFBfBrvH2V9onoy1xlL3O57I1J8/+L7GEJrK2zr5cgPvS3uQwZM9SPGzsfT73ysV4UUrJd602YJX46KbSuJ5j6u
ObkPppCcxRZy4wuIuLJtX75FLb3cyk6Rdtr2YrOTwi6RmbVYK1qjuoXAlsggNnPisXgdWmARIacxWQXjUSwxyQMuppOwAelCWmHFyWkURNH19lJw7isxNbZo6b6xjhHP
1UgSbBANq1I5LpQUFsDmHNRVclfbArlsm2JFHh4aUON4ySeDqWbxMedA4/1lURaZwAnhS9e4yfA/ecGkTnwtcYIJfDVEo+7Z5/B+lDMpQ7hJVMTIEv9nsc874lF2KdjA
QGO/TCA4WafH60OJmscU2JjOEuBj9H527cVvjOnTNrq9Bg+8aKue9zQCB4gZ86eAvibmQeL0hwifjjR2aNWzJz+r9esPW31QZRJSvwlbT0kZY2h353Bk3YdT0zhlWkhh
7mboEgjOyXeZIG/wMpQuG8zgmzG67ohgYI5fr/g0CGdJVMTIEv9nsc874lF2KdjAvWuflrsGifuls1xVzS9yuEg3ZTPo/GDb6GC2Tm7XjWw3vdJCNNf2eIr6Je+nHAfP
280nS3hWBZCdOwNMO6NLBe4i3IOgyPGh6IRollGPDpEGbWA4nH0QJ2urx2L+EnQRTNRs9sZQQ8JaSXBa3ar4MXCB4UlDpdMdRPWcXUy0bleSN+uUxOssSsbeJYJ+FM0p
L00+VoF00p1m4QPt4caPxvX2UnDuKzE1tmjpvrGOEc/8WuuaRFTxMjMQ+6GQ5iwPfnC79jW+QRvErUDew1vqfjSlETbBIdwV/VBglBvCX5h9YbXSO+PBxWcDP/niyz/w
280nS3hWBZCdOwNMO6NLBYkF9j58Km6llVofyEEBLFmCCXw1RKPu2efwfpQzKUO4280nS3hWBZCdOwNMO6NLBS1+6akvhS72kB7UtXPAlBhflJBNir4FVRiH4i0vRnBs
VB8e2K9tb3XyNaGbGWJCCf37+aOlW5xDmR8hflri3PgiWKh+4/gmQGm0y5FU8KatHD1CKb/YQYeorHkoA/KbCKTWniUMsslvH9BQHIr1L/EKd1O26NIE42P0dpYMSMVO
+pwtS6w5SNDK54TverUTvAfttJlmpuvwLzjnzf5sLtGBkXrO9qKx09dke64T8wy+72vnXapoeiGMtDN1I3R6Q5tJEM4KoB7c/gxrn0VfHEpBLIbatutxP0VgWLgNOgPM
mZ6ReY14pkWwdTIORCU8QSbg01VSwIr0bICzDu1Iu27WimvusHDbyMQ41+dZJGia01LnFluPjQriFnxrkHZQ9EYRryYDAmrMm/WbF7b0lmwJm8zxMW4UKQIE0Yv0qo8g
05VjElnj/f+dIiB5pOSgdVQfHtivbW918jWhmxliQgkXcu1ku6lQOIETrZZ1IX0PI1J8/+L7GEJrK2zr5cgPvfzF9rwufWaZBQOGyMy0CdXjdC+ap9Vgprf8sAfiA25q
qKr5dNaLOs41AvYFbz2ma9OZrTjTXjjj+CPAU9cPFuzbzSdLeFYFkJ07A0w7o0sFmHK2y1QOzhVNTcfyJEXZfbF4HVpgESGnMVkF41EsMclzlXvCy7MJVl8qMVyAYKSm
1WiiHmKRGLBaxq421KPMrhljaHfncGTdh1PTOGVaSGGg3esjFs+gog2w7/rBbVePP6v16w9bfVBlElK/CVtPSRljaHfncGTdh1PTOGVaSGEsej8XZLelYtIkkyOOTo8F
DiZwihgJYNtTpJSdgA/wZ2lpXbyTaTNJaBoKFo7MbcwbDMb8GnoAne2//80qLEKuejf+mRt+vYb0P3Ur6tj/wj8+pD/vXeHmSSfkiLGc6k9UHx7Yr21vdfI1oZsZYkIJ
Kp3npejnLD41ibKG3p7WTQhp+03e655OtqDrsYO3Jy6k1p4lDLLJbx/QUByK9S/xJhDVvr4DAwHCLuVoeacujNviQpXtprMfL1fvUaByRdhTxAiO8QVm+SmWHDr0x0/g
vkUtvdzKTpF22vZis5PCLjAarG1kTQjK3eqsDSjKOoykVZJbstPKCIog6ADO/T2/MsoO3wfXyrMxDiRpA/b3b41h6zQ0cT0f0x6V3E0sRLMtAR+9psMefgVhxn8tRXHr
cnDxWPaILTh8fM/7FSib6YI4MObJhhT+e0T9PeTuQQdpaV28k2kzSWgaChaOzG3MusT7D22e3HkJv//SO4QKI0cqx8jSfYn+ic9Zys57YUU11bUaWzXWWUim/QYr/Jli
zRDOA3k3MDV3I9PV8650vpzsQQ4lMeYgkJkeSZgbTZ/+iHbkx90hwuQ3TajI4Zn2QSyG2rbrcT9FYFi4DToDzGGfB9DfsBb15Hk1hWFFQxbr2EctEPIgGkscaKjmIjvn
yFsTygNU349lzX4Hm0k1MlL2y9Tzrsr/OpNV2B9vyrq+RS293MpOkXba9mKzk8IuUK5ojc9tAgumRwQPhjapFlPECI7xBWb5KZYcOvTHT+C+RS293MpOkXba9mKzk8Iu
CiRzX4ifWwqWgLeRe3q/2NdfJyrwf1Ottegc9XmcjCkH7bSZZqbr8C84583+bC7RhH1NmoBaqirsETsV0OKFtiWOAv7B8s/LBBZDPhCMDPPP3BMW10qLA2J5wAt4y2aZ
MsoO3wfXyrMxDiRpA/b3b+jMmOb6GXqSuXRndcww2fPjXwtcdEuvKhuL2lgwKtXN1opr7rBw28jEONfnWSRomqPFL+FaUfPZ+60HNcz2UwO3i4Ig2PL0VqDgQdS7yMrh
ivQDyagDc706yuJPXr6NeSa8qayw7H1r43fSDmjLEagXI2F/j59yR4t7ltqTMLZBDKcTDiGhNsnLhVo06n6Yza3hTU8nV5EqbIYJIbqx8jO8IwmG0eIjcKlw2WuikbHa
nHQPTFnlWAPAgfTYzL+Kzzo9AXChgxm+xg5inbOt/1V1siXEpye7BR39rSreNMDVbSDhN5Q8jaPKJVrJS3woLfNsOBGl+w30PbDnxp3j+4ric9fm+UAg8fl+7/o22bSG
bycgxdeeVqercBcNqAFJ52TSyc8RFkMUhaiRHAnFlrZY08x2omlJS1xXS5KLv9kNQSyG2rbrcT9FYFi4DToDzNpxWec5AvWeZxkeOrdaMP5MzIoxyxqhw5h35CoCADUF
P6v16w9bfVBlElK/CVtPSY93GlelYSL5HhVUeE1xnaaQ0V2TjN2U2DHVmDNxLjLzvmb1ladDvcyEq4a5t03B0HZiKApPP+EeM/iSMgSJQlE3Qp0FtJDYtsCS8o2wG7RT
+aZsXXZrxlMVI2CLxpf0thUrd4Rnl8wjOL9thY6XoKkj4ojuqOJu+kDBIlwf5rJsB+20mWam6/AvOOfN/mwu0cxR7hiLNp47ub3/WS/Gfh0/PqQ/713h5kkn5IixnOpP
VB8e2K9tb3XyNaGbGWJCCf37+aOlW5xDmR8hflri3PhonshG37pJG3Y8AgZUjnX+PRxo4I7iEBFn+KMJcUJUi2dIJnJrYyuzr+NhL/u573Eyxc9U+/KSp7rDKGnGxKtm
pNaeJQyyyW8f0FAcivUv8SYQ1b6+AwMBwi7laHmnLoynphJRwnK06j6eR0SBJ2uMumKaxB3Vkt16P3SUsQ+oHQMuppOwAelCWmHFyWkURNH19lJw7isxNbZo6b6xjhHP
c7E9lqLvRmrItVzqrrxV8x5jmAgMVoP3pRnURagwITs/PqQ/713h5kkn5IixnOpPVB8e2K9tb3XyNaGbGWJCCeNb6Lk+8rCZ7WFDw89qyxXDDGgUQVvXxZJzTIA0E7ON
odj21CDpAptH/aJGsU5ecJDeokS0xyfpFA777A519NMmvKmssOx9a+N30g5oyxGoFyNhf4+fckeLe5bakzC2QZfWaY8wXFXtOkcWtOeiRNOyDeGtse34TQy8Q6qYaIpZ
O+43zAOjMywxKbJ8K4J2ab5FLb3cyk6Rdtr2YrOTwi4KJHNfiJ9bCpaAt5F7er/Y96e2ZpB7TuHcJXhEdzYFl3cR153sF1LSjf5LId8D6EUcPUIpv9hBh6iseSgD8psI
pNaeJQyyyW8f0FAcivUv8YXBjl/PzvoR3yvUzNd2EIF11MWoC9QepuAGacisDAMmAy6mk7AB6UJaYcXJaRRE0fX2UnDuKzE1tmjpvrGOEc9NbkZk3Vp47RAVc1rgjxHQ
bofkDizG/lmlmn4DuyqbkqgIhbAcDIAbaGkZt2LREVPyHz2kS6G7LoHFKLjHNyE1pNaeJQyyyW8f0FAcivUv8XaLNgrSyzZKxslH09KH9HkM605Ce32ZSXhOiyuFVkcO
U4rwrnFUipK5eBCTHjsU/EFWxV/IzUUS9TFuZp5TyeN9vWZ4zzMG3cl0t4VLP1XWMsoO3wfXyrMxDiRpA/b3bx6FhBpXCFByoI72IeJiL3cl6YhGoXBz7i8VUYG3VgQo
zbHAFgrIXaPEmKvPIJ6kxtaKa+6wcNvIxDjX51kkaJrsJcKkgyxin2O5Jrqz/ypc40/f0OHYDQ/DcRgoIDaCkbS3/GKlDJ0xkK9jC1EYO8tS0KozC6YS8+TNnxXrXurQ
gbjx1FJxyyawsrVS85wLh4hlyPMAWs3PxOQeQJOj7/PzbDgRpfsN9D2w58ad4/uK6C20/69YW2nx4GGHCncia+iDUHM7covfhX8R/sQiZfE/PqQ/713h5kkn5IixnOpP
37vlYxtdCeEOwhog7srFsZ7uPGj7H/ne2yCYxgqvy1/abjq2cJzn/2LQY8rf0WsHwYmXbjYo0MIpxRAE1XWNftgm4DFgfxxqviw7uIgpjF8rQgQz/Hhn8CaaJFoibOeF
OeQczoyQFmWbfE1aF8BLl3/vYJQMm0Fuzb+cy6CHDx3gfvDPIL44o4Fd03QNnc2bfLKc6sElkKtAIsLlJsqgMtaKa+6wcNvIxDjX51kkaJo8ChtrK7FtzN4wEPeUfDGy
v0vNSMGK6PHs/dX5FjtPihUrd4Rnl8wjOL9thY6XoKnD/JVh5V2xGuG2HCHbD89fE+SUl7h/k84NB1ynRHJU0zMdqnTHEoS5ecYZtvj72r1HLvQ2de8qJj2zMu2VcSC/
B+20mWam6/AvOOfN/mwu0V6MB7RrkBSh0uLNKkgpXdhkWSw9lHZYU+RTEV5E7w/KxyQ41SLt7x+3raGn6w84tdKcRz49trRooAAcgWslHwoKD7GdbzcSltr3aF/e/s0o
MR/aBMmyQW5O0lLFLqVK9mJu4OJ43r/pgsYnaHd3zJIhZBLs/smAEBo/o1E9ekiR7rJ1277mcl27XPNtbYxQx5KRRAB7wMSHGSULJGxv9FaM0uGyohsqBWKw4es0BJIi
nRu+6k9KS/9uQT10PQ6gcu2Uy7QCaM14v+axNvRYdadFha3BqO/K6nU5OevzxoBQjV2ZslN2fnEWoOW0oo4Errp8jBxM2v1FYDb+KT4N42F6tox6npPn6JB41lj0ozK7
d4CuP8AoahZYiVxhyKGxA2jIIpFvWYVZacbpx8vx8ce54mUrNogou2XnrEaCECRUm7OUpyqr9qjffPe27Ox6ApQHQaYbbvQf1Pt9avxEeOwHF9R+VqtndpOEyXql+XFG
2g+tGKSpDNkJVIzkZHuRyKgIhbAcDIAbaGkZt2LREVNCIFCO/cnEA84w+RB7GNegbCu59zn60po4R62ZOh5ZC+6O5Uv8+UkeI9fToSEJBXUucdKVh4ipgxv95DZ4jhP6
s03f5MYVeA5+kG9WJ1A6Ut1ennDBQyr8w1swTXHoGF4zDFK3oCfMLc62Tc+xRwtRG0xozCj4UNRgCKgHERm+inTJjLFJwmbiMOUY7oo10Nq2Ce9AJ9S+Q3pIy2nvyaxw
NtBu7+/YsDdx4H3xjoiWW+zHRb72D4Z3UnP2s9A6DIdH+wdJqpifnnOOFz6d/GaFccNGD9HMG1SLUnWdioDfB9yzlAXaLTwWJ8PzAsjRPH0oCyA6rbNwJ8vsTjND3aVx
7RzooaHyfF97YvjIDpihUtyzlAXaLTwWJ8PzAsjRPH0ldzO5UQImPUBEbfCiZtfelCHMWJqJm+g/+OGcXAbvxNyzlAXaLTwWJ8PzAsjRPH3rYFREvwEDP+cwSlNhSIIU
qNUD8n5TxAREYxACFZ0astyzlAXaLTwWJ8PzAsjRPH3S0Xu/7uFVnxyLNGiu3W+t+fVzGtpBBz9AnQvJZK43i9yzlAXaLTwWJ8PzAsjRPH0B1fL+EaAcnBGF8Lz7vT0n
RWDXWawh2Pl4kNKjHb8Z/lbWFbJMWQjuZ22pOl3tr/nzLJup3x/2Z+xjdyymrXEE82w4EaX7DfQ9sOfGneP7itGIrIVGaqWCc6gp9RGq/RYtCTYKkEcZ+2oY2hGo+1ot
IAIBywkfLXkVipNm/PHgyLQmaqVkUnGHp/0Bda8vL301Fseu7gT70q1Qm6EK7K9lqfhtxR9aVwI30vQ/mIF4Ke0lj0NE1doS9OCdV7dLD6r4NKl+rHeF6jVL6Xw8rMzt
dS+H7O14Wpc11dObnxWBs2bsMd/bw3IjyL9vmLLGPR6gSLU++qFcXmL5Y7fFlpSYtxvFv0NomDNMbGYcduuh6Z2DuYNdd6CORZMfwyL7eceLXVZHhtiT+/pBCzv3nfXC
nicTaYBqJ2SgQovHWIXURxNNwpu5In1wNPj1bx8tzVR8kYLY4DyAFQj2HYOhA+33wgQpyMROFJZW1b5oZHyWGjIi8dTOTkS3zzCJCQV+kuRTeLbEXbgWm3CLkJYXA4be
ThsG2KhlkWHvmLYjsh4wO2yrB1A8u42FK1SotkJ1mMVTeLbEXbgWm3CLkJYXA4be8Ix8pefP2AoRXOcVm1yWTBlGj5GKmqtmy0t1AQTT0YVTeLbEXbgWm3CLkJYXA4be
qTD747MubujxEsHvXUATvRAScVooanjeYHK56xP7PvZTeLbEXbgWm3CLkJYXA4beV+6yxIwZ5AcJd0yFRkuv7kKAcpBTcuDVw+idg5daWhNTeLbEXbgWm3CLkJYXA4be
jFeZeIBkkGn4uQ7VhkP7nWrnJGZQ88O2IlF/aKFulWM8ZAL69m+Tc4+LwxtOpx8FCZvM8TFuFCkCBNGL9KqPIKNhdfR5Fp4Q5c+GCT4xdBX7Jlc7o5UCfwzwY8xvhQnt
saK3iKrZZbd3KnILDHc9KTuykqx0gfcICiyuzaJkxKTvUptwsnXPU20tcFeKYlikZIjTOOfXNI52/h5MG3DGmszLFhvJEoiy/sqcNN9H7pLIPjCIEgbr7SsclOLNGPnD
GYP+g3+xRfxdYhg2YaamGi9DgB0M02N3O9zxppGqWw3Lp8VdIhBWAFNTpV7htjNWM7GQJpwRZgh4SWeCrfVKtBDv4cygclaijBu6qAP3iL4/4wnz2txHFZOEVQotSFd8
3KqHwPnVMICTpYbOv16OovsmVzujlQJ/DPBjzG+FCe3+NeEqU+zDkG6nT2FTHfU3unKbYbGcspRE+ZjdAM8bTvsmVzujlQJ/DPBjzG+FCe29H4m5kor5l205bKob8gxC
HjaJ/tyUJeXnN0ocCmf4cPsmVzujlQJ/DPBjzG+FCe2dDfRwgIMjxhnwUaOOauKu5/KyfBvRGn13U753Up7Ji/smVzujlQJ/DPBjzG+FCe3q2altj45saCISwMRW2gUd
vYk90F903IP79HT5ajrsEvsmVzujlQJ/DPBjzG+FCe2Er3dJNQoyeMVuxiMYcXHKYu1ofrgjmCuatET5fTOz4qQ4MzIv9e7fNFzEV65MEoxDlCBlV38s4T6SN1F1R332
qzsM5KOPZqL2GyJNnVBAhOkZAvOcMbFOORCMpsg2sMDGSJQvx1JaOZzKmlkEYxpWVIi1P0Bkptg52e7nJVXHMbPqzge+g22Bp+dJaQJvBsDz9+N1IQiYxFk+00ZOkx7J
X8Q9kEuxJoWpHJ12QDsQh6ieKiXUHoQ0whcajYEkEgbVaQgrTd4eSR0QL7oZUad1juYHq5VC+sfnfrVLbaFfcj8+pD/vXeHmSSfkiLGc6k+6nyRHPNkJ18QrKqjuoCGt
+72o7WfXIOJWp550QwYjq9XGiwypsKvBfsYyyOxolKCu7pfvXxyBj0KPLmN7P2KLzOgUErPd7ZUux8aJ6sk55CXAoGyKbJwYleWX7W0LL4yXt3V9yTVaU5UozyMJM0kK
mWIZdoaIglWWIeZsDodWVZmkWSdpNlLErY6M3XIlfLH1nPTdhFXT/ZZb3cjyxXMD7yo7sR+Dybc2G8tOs1DEjaRD3rxE0dV9wuPVssHpqkArna0c3DSZuh3Hfnd/Sr2H
Nb1vmKnI5FJiuONNh3s/kGHdbsjkgYa98KjjLuA8dqoixuLas4nue4k6qL7MuXnFNb1vmKnI5FJiuONNh3s/kFjWIpfB0jJycLQlP01e/dCwINjE0hCHxBpzjtMh0tT9
Nb1vmKnI5FJiuONNh3s/kHxo8/W6M6L2huqZUG0fkmA93Nswo6orf58nhv/sgWiCNb1vmKnI5FJiuONNh3s/kKzoxZSFVtrc+DAK18x7UXu6HNvDjYbAJhjJyX22cyTg
Nb1vmKnI5FJiuONNh3s/kAuyC0nOyVGpCmSDZtzMrPBnKMD5jCz+1k+UA/BFpqudtz/MSUExFCo3YSxm1/EC4BNNwpu5In1wNPj1bx8tzVRyNW4ATycUj2kGYveDO3yS
sgIK4tEKRklouhJHvhrmxCPKDKpZmtxsU8vN5B6cQ0TUfvTWZCtaW+JkeFAyJuHhpYAU40a2mfknRk5FEzg54HMFIYYerQG3v0XlnStsaTmGlA4cv080jvJS31Yf4/d0
ba31JGXhEh4Mx4+Bj8AbUbewMS4KDHx5V45y+GPsCipN9rW/AZ7YcstsSL0RVNbIxC2dIh4APZfR0JddIg52PMHamvb51TCHM9hqqTH+GSioXj78Vt2hPyqqgK+iiHaa
FnukJl0A4A62i/nSw8Jr7zmolU/zG8j25i2du4QjfWLfOS4pyoFH2EVKH6Okde3LNB3fg5w3LudQZi9f+NjDxTmolU/zG8j25i2du4QjfWIkyK2SUFC0ym2HGrsCbnYF
rPRf7zxZfsOmrqduxMt/HjmolU/zG8j25i2du4QjfWJhtVZpdEaiRnlNnCTkoKLulOu5y7hQ+cm+rMZofAliIjmolU/zG8j25i2du4QjfWLd2xJcAPj2AqCW7J6ebxCo
EyysffpYALCnqAo5AX7a0jmolU/zG8j25i2du4QjfWI4Zz/BQJI+iiRbKXAGtOud5t0BmhA/19Aibqygp/TIs0F2HR2yqRd2A3AcRZkDAEkHHk/ynKRr71LABjKbi9ve
yWlaUNmiiAyz0lPy3BtIohSZaybawd4vkoWZsIWLiXvQ9Em4goepiMsnCZlJZl9Xy5w9XdMNu3Jak1E86Z2Vdz3B22G6nnHz4c5VeqKl9qfXtpNtliouSSkh3/JVp8Kr
CIvGrCbGwVxgADLaUiY7t3RVu1DqJo99cYThzb/wnuilKdOjauwGsPaPeOp8RIpodiSaBKLeh0buzUVbI/vx1jGz/+Ggnzm/qF7Q5dI/3QEi+U1/Vk6WMICnK/eXhgvc
FcGwTDDrawtgkehkCfxPRcE46Mx7+TKxHySeS1PIJw220xbNGIzJP/sRi3nPdyxWS3zOS+jhHvyb+Aa6rMKc5G7H7NLun9HQU49AnzpZJ3sUMA7sMe2OQekSpwnQwHFc
5wi9bTE+8+lq/jkWCdAby1A8wEcKE+mMBIJ+CATpdlIqCWoa3nogjwy5269QqWanun46cpn2PNsnmX9/MHF3lAmbzPExbhQpAgTRi/SqjyC2JIl4KMts7JrSQzyW0Txz
SEiMK5J/opqig/tBQ7CtNioJahreeiCPDLnbr1CpZqeMjW7BPgVxv0+RwPJMgiBjL0BrifRthjkhwcSYRlkHb29IXBDbfdgXnCSuCWUEie21l0G3J+2IKlNEOCRgBmWD
TErX1nXyNpLpi3oNUJM9ilCQn4DAgTOd55QuaQD1oGCE6YAZwfC1+JILDqbOegZJTNRs9sZQQ8JaSXBa3ar4MT6SMC0ZSK1ABVT+re4XKVIDLqaTsAHpQlphxclpFETR
YyyuaAR/BKy34Lj07ulbpQtpMIMgZIaNvZcAAgjJjNwwdrgnKKeeDH7FpOXepJ0D4la6H4ICiXJooSgb/6dnNvX2UnDuKzE1tmjpvrGOEc/VSBJsEA2rUjkulBQWwOYc
4vQ11WDKbxap7tZbG+MHA0R4X7kDEIbf0Xvp3nKvk0a8NNArBwe9C0A2xGbTtvdhQtiphK+CzxdNeskmnoeuH7olYxZSn8wPeDg2VgzjnQlUHx7Yr21vdfI1oZsZYkIJ
WGZ7POj+s9vqVJGenlClW7SRJ+hK7AKyBz44F0D2GM2hxAFjfu2C9nKAbgR89V48WnCvfjIq8KfXoYBINNCbEL20JLyFzXQq4YeGK7XoZeuny0JAJB6CI5o2HCiDNQKq
9fZScO4rMTW2aOm+sY4Rz3OxPZai70ZqyLVc6q68VfMZooZIV/wWel+gpQqC04mInfQA6+qNU7rGv2s/Hmbaxr5FLb3cyk6Rdtr2YrOTwi4KJHNfiJ9bCpaAt5F7er/Y
HhzAL2X29ToMq56fXNQCEhotccfsdKhpnNnel5ePxaeV8trzCc6vLxV/IjF/HA3zBnvUM6q1qOT5E9EFiUhlR8fJJlNip3Z03IG7FvkHlC0H7bSZZqbr8C84583+bC7R
KDRx7JxP8q6BDcVBzLKgAkOdANPLqN6+DMYujB0ob6x73bPvvrIEdgvMOAXfI6x458GQi0JXTX7ZqSvNlpq7neQXKcuSLEwZRMKg678x0Hc+QdYZXDNItl+EK+IkTAk9
GQ5YWqnEiIsepVPYoWbfaZqJqyZMhsWUCFGxO4XNOGjBRPCFsvnlIcIQb461TURCG9vl15TIuCdga3JpSNFFhdmnzO0JeJ3WlpG6DaI5liPiGVxY/kzNIP8hvG6Q6rNr
AMH48TyqFxlAQJNLREwBxi3uQwZM9SPGzsfT73ysV4XmnhW3CcwKrx+D4nKlWcuNk8V77BuBaAXweoRCX6dnbUQDd+Dr6qpbSuXO0fTiUTXzbDgRpfsN9D2w58ad4/uK
uU1O1hvLRlBOPD4GFM9GcRn/wxWElJHHjYq7i9XTW8e/Zynk4eEH40eiiYpBmmb5fb1meM8zBt3JdLeFSz9V1i3uQwZM9SPGzsfT73ysV4XmnhW3CcwKrx+D4nKlWcuN
xSnWmw8SqfdojSYPzGyP+AmbzPExbhQpAgTRi/SqjyCO2ZTe2ZGB16Rcv+0Hk2vJV31Nw2rrCMSC2JUKblubLJ/rigpR7eE315oBXvZH8vIRZ/5zz0Dnt+XYeEgc1lAs
VbcC6Tn8V24xFIMZ8VT/GQ1rEjat2MhXCEvWr58k0JNgqDNVhtYGo+9NpKrb+GwbWDcHSCAYMHvALeH6nO1/eaTQ/pcUeRgwGH7m+0IpBnj6TKnsRDdUgZETqEJiDdrM
laVSsdyJi16WXcKZbNgid/wr+TA1/HGALKXr17qTuLFrSRE9uOAq5udFwJtgFIeh0KjkwqVuhWVEhY8KxqDMAGBA1Nx/M+xlnDQLCdokPJIFAeo2Jj++TUJRHs53JrVY
/oh25MfdIcLkN02oyOGZ9mtJET244Crm50XAm2AUh6HQqOTCpW6FZUSFjwrGoMwAK+IFk8uUj9CGdgRKgc75ZKTWniUMsslvH9BQHIr1L/H+IrzuBFVkugRmRpU/gXa2
RUVp4dcA/Y0fdoDZ5Dp69jrq7CGOCNS35wEtOggBWq/Tma0401444/gjwFPXDxbsC4UraSjHafpcQlHCMykFzjgOMLTuWlFsGZ29c9wT9OWt4U1PJ1eRKmyGCSG6sfIz
fBiuKKxARlTaKXFzQvSG8tufsH9AMjHBxXizj+gyn+eqZgf1Sru0vgMtJIeqEpMbde2+DjsHQBgazTzRq5kaMAU5rHA6jTipFiK9ZkUHA0Z05NmdZBmm6Lzfk26ZNkOk
G0L9rKq0ORdYZu9vw2pcHlpkJoYaWzJX3NM8piB/6zHP6C1vSKfCbxj6GMSTj/KyObkPppCcxRZy4wuIuLJtX1ckXuxLcCqmo+ANz2t69gm/ekfy6LSld+shoG/iPJTQ
bvVRKOCo4fpic66v6ObayKt+JSwRORMjo4ZlHLxhcBVFD0HxhLEOS0NIC/hrFuUSzCrOmMP9PtPMSsvDb4hj/gU5rHA6jTipFiK9ZkUHA0Z05NmdZBmm6Lzfk26ZNkOk
G0L9rKq0ORdYZu9vw2pcHul1Nt8JQb3IjEBCkziiX/6n7G2L1+gBl8Fn5NwW8MjaJryprLDsfWvjd9IOaMsRqK87xwTmFMFQqMLH3BoSJ47khMh63po1IBJJLrNR3ekG
Q2Ra9WfjO+yIIf2sbM0UbfX2UnDuKzE1tmjpvrGOEc9NbkZk3Vp47RAVc1rgjxHQG0OZnk1PEbN3P3LCLi9FnzXQVKB58yu0kZN6j9QSYP3zbDgRpfsN9D2w58ad4/uK
vK7Cbt+Gi+yt9ooki/gaISviBZPLlI/QhnYESoHO+WSk1p4lDLLJbx/QUByK9S/xxz9MAn78i0+uS3r7GOFpTfDcihht22Sz0lPxR9ydf8ImvKmssOx9a+N30g5oyxGo
FyNhf4+fckeLe5bakzC2QfRZ5UCN+9kN92Exip/BseLzbDgRpfsN9D2w58ad4/uKvK7Cbt+Gi+yt9ooki/gaITCArGDrXND+gHn8go+hNAjWimvusHDbyMQ41+dZJGia
VeaoZw2RsJSqJYaNYNA0px/0CHNcxa3O+rR5qDOh8Iopd3LXtg6zBKY+w08UgeDlpA5rlaC1sFOTZ6DPVgB2sslUWaimnzh1CWXiqpYCmJ0/q/XrD1t9UGUSUr8JW09J
zYe21piIB2Sv4L+vEC4IUznncKMfyYBqGLnQcO7UITbzbDgRpfsN9D2w58ad4/uKE2jAl2KbqYJcHYVkWCpkduhF5hLqW61fzHj9eKYDMqWGGubq3H9F7b+qkLChK80b
X7aLw9jhUcNJ61wZcmMaWfMn2isDdIO8Wg/vvoueOEQmvKmssOx9a+N30g5oyxGoqJZQ31/O0KyVp8X9pZuqz8u21JTY2QF7PRKRGmTDTWGrwwYqSV5ywX1G03Zudv2z
1opr7rBw28jEONfnWSRomrdadAlmmYa35Pw0eWnTdgiTP7fDRVcJIy73+ezVr+jLTNRs9sZQQ8JaSXBa3ar4MRTfxPecXOFt1mQqS3Uniu23WnQJZpmGt+T8NHlp03YI
fTO+u4w4Xgy/wa0JEqr3FwceT/KcpGvvUsAGMpuL294cyZcG2G4P5kv6ZEn4fQSEtmxB29c43cpukrl2PpxJuil3cte2DrMEpj7DTxSB4OWkDmuVoLWwU5NnoM9WAHay
WMW7C0VBGZR1yr5kTaW1WGmoEoSp8R/pwOYK1bJShrZYjGYTrfqLMKDsMKwP7Cw3DbYsu7C9SF70UGqlhG7LBeYDeNp5u3If2/KQSzgeR5S1l0G3J+2IKlNEOCRgBmWD
MXxKN/2cRm4KfgZKi/Sd1lIVpRyHzl3vGOnIdWoh5VtcdXNkdWcDPAk6PVTxHCDRy1jPIUmezd9DZe8Y5m6aSJoQfAOdn96zE5ilZf22c5qrD2EZ5b1Qfxl/AonQ03XV
mdmrFZzGccbqdNXNEc0QK2/WUoMdI8CDkzmFhti+E27XlmJzEgSBYumT4ZpFnEhKg5JZ3VKRJj23EGkjcKL7gO9z0Fkv1yM6X9vd1tnMQtGbnMoNAodGABpp0FYbuHZB
+w8RLP+ui9m35lOkVWOpxnrkOlCLFbx0FrFqnRcuWVhoY9EPHP3TP8Dzyshya/i6wULQDOP8/kUB5R3wz2I1cKUKey8Hxt/3RNH0yFLFdjdcAuUM01lxVo/JvmldvAKy
vIAmVtoIQ13bGKODxpGLOhndIu+OxkpCs5bbyCeO+h3Apva2zJyZfH9FFMjS/MYYlbmvIi3mhvy2vtqvpgapYyfJwCteUJiUFB6IcCwJW/CCN1ro9TMW6EryAybloWE3
AE5xKUvB2zCtWyoS3DmJXaXRkHDi+q/dDaMwURmAQ7TW+jU51eNf5DQxKf67RVZqm5zKDQKHRgAaadBWG7h2QTg0Ad8bHTH0O9V5v3Ii0s1ZjpMOMSTea5q7z/3V9luO
m5zKDQKHRgAaadBWG7h2QdtMX6rh6KBJoY6voQDXu8JNnkN3cRs1ZIttgB112KuH7FijRTteRGxpxlmxx+1ptmM0GrLNItTGRwV7bq4uemM6TK2UmIj0C8gRl/n2miri
PurMoCztlr9qgwTA7okVASfJwCteUJiUFB6IcCwJW/AkOoxuHJA1hR4Zk8a8600pSG2+txuyWmHYlCUJKIAmv9VjktKNFMTRVTCLTnvlI6jlKnDs2fCcIv4aeXtkrGeW
vWArRUsaIQTyt6HH1y1m2iZP3FTxAhsPQcHUu9dxPpZYI4UWcL116GkSBuhdHTYHP6wc1BJGhPu0W1Ec+KWb/VvkTPSt0p/FInGtDFUXLu9cAuUM01lxVo/JvmldvAKy
vIAmVtoIQ13bGKODxpGLOn7KPofeI7m+a/Bmumb8bP0b3MtS9qIedjbjdYxCBj/THaFK4dbm8HpFbTsHc4pM7Whj0Q8c/dM/wPPKyHJr+LpQN/PynUYQCimryhUAh6Lp
w7LZgOFdjs2S3gMSfhkEUl8ety5odskffEx8COird8JToeqEIRC4/7ycPkAq/OqKTZ5Dd3EbNWSLbYAdddirh3EHFErppmd2Lz2lv+fbEYivhZRuA1PEuBomdKOGdjDG
1WOS0o0UxNFVMItOe+UjqOUqcOzZ8Jwi/hp5e2SsZ5a9YCtFSxohBPK3ocfXLWbaJk/cVPECGw9BwdS713E+lmKotDnvmTQmqCETEwnsGI5cAuUM01lxVo/JvmldvAKy
9G7XvF35GjErYhNDz5Ohgb1gK0VLGiEE8rehx9ctZtqEM0AiQl4hrFby19oUN2dg6rdiCytPbptOJaqRMG0FMSfJwCteUJiUFB6IcCwJW/D2xchLpXha9IS1ZDB1w9VG
sc/1OXOHR1EDxDayD8CkMI3iPphrYl0fidWtVjKz02ElE7BeB/w2qLek8i355O2XJ8nAK15QmJQUHohwLAlb8M5qrqxX8M1tO00SeQX42BhoY9EPHP3TP8Dzyshya/i6
R7cZJ/iOtlpIrb66Fj2WE0zr7MUsp1op7iBdjTbo3sdxUpBKfaN+O5jlV9qg2V1fvUJtkNaSdFIv5POtiXDY/oXdpGqHOoNlnsGGUGAp7mzRFw+Q42uZ8ytx4IbG0ZOQ
b9ZSgx0jwIOTOYWG2L4Tbm6C4X4mzphbxUizRg7nfihwKDRYjNirXWLwT6mZ5p0XwKb2tsycmXx/RRTI0vzGGGYmYB0z5dqydqI27Fe0vvXiqZQZvHcqEYCk87jlmQfg
m5zKDQKHRgAaadBWG7h2QTd9+ykY83thG6CTCcgYo5/4pua6Odp/becoIAdOL3291WOS0o0UxNFVMItOe+UjqEC33DcFlcqpUzxSSseqXDnG96H0sa5TH23fKCcvPqFx
m5zKDQKHRgAaadBWG7h2Qbtuz42U1AXkK8qVYyP7lh3FbRKoXJ+94P3/vbN4aivOXALlDNNZcVaPyb5pXbwCsrLhoGOLpatml9mCgyzNYSN9O+UYPCwMew4psN/fx8qe
XALlDNNZcVaPyb5pXbwCsrLhoGOLpatml9mCgyzNYSM9V29U5UoTIQGRaHhUfQTwnXo95StI6rHAk24LA0vVNFHxQVN7WuZFmQcNCEaT3iJmaL5shwKiUv3ag3eIrkjL
Qhd7/5kVrjCWPoJACkomjpucyg0Ch0YAGmnQVhu4dkG7bs+NlNQF5CvKlWMj+5YdeyEBqAIJSbfyqXdqGCVdwU3fU3B+6mUtLmTXx4iHcxl3T7GFBhyxNcRYGKUCQz46
GNbLhFAChgACEX4uy3VbfE2eQ3dxGzVki22AHXXYq4c6mHABMu1oDkLQSgigrVX0sMKIyL3aDaRUECYumGybW8QLl/H7dq+gR8Dzgb1ly5/S15y4dWbUQPIt4bNC2dHB
fgy+udCwAxFpwmPGLuYWQjkuGhIPwMTqo7Pva39Ji7WN4j6Ya2JdH4nVrVYys9NhIqeLZk7r7eua92aXU5JOxu7ZF9NrfVzYl9doXF0P5w5N31NwfuplLS5k18eIh3MZ
d0+xhQYcsTXEWBilAkM+OhVJX/xqOKcp5j6rD1UsabZNnkN3cRs1ZIttgB112KuHOphwATLtaA5C0EoIoK1V9NPjkXCEbjC4gNEk8MKGCrSV2appuvYpZCi9xSBA2dnk
4qmUGbx3KhGApPO45ZkH4Jucyg0Ch0YAGmnQVhu4dkEMXLXkqv+d+M305iasIwSS5nA2FVfxPUuowlXvrYkYXxvcy1L2oh52NuN1jEIGP9PDThk0HSbbuy/SuJkQkbxp
Ci/y6fyILvLYx7Tj72E8KLMxvIL9R8kq71OuGA5B1GfQ+BBG1S8pM2jYALWcT3G7XALlDNNZcVaPyb5pXbwCsrLhoGOLpatml9mCgyzNYSP35QUxNG5ytiyaFSzz/0qy
99jsTlvZt5R+Jvxiwvr5271gK0VLGiEE8rehx9ctZtqbVrYkBIkFD4X62YA6Pf7Cr6GYMIjTzsj8w0EdAgupCz+BQPH/w+RW5XTOhCpS0+w1jO7yAou0B4SAI7MPKx6H
A3YetUVcRYbuOkhPjxRyDHe/unM/Rl2YKkFLqHiJTxE3hVPzDvF9uUMoIU9VG14qn1qp1AczyU/hfcGKotdzYRvcy1L2oh52NuN1jEIGP9PDThk0HSbbuy/SuJkQkbxp
2e41Q2OMUT8F7Z7UZCqJcTJvgVPlt7nK6CdOKLtmVgxN31NwfuplLS5k18eIh3MZd0+xhQYcsTXEWBilAkM+OheucbLKjkmrJI9ei17oqFyl+Voc3gfHKbxpvFaHmC9x
8ytkf2e7k4C1qfq7qLXcT43iPphrYl0fidWtVjKz02GE5h1nqwZbfc8QzZDh4OM+GfbENJ91F8wW1HtgNt1vw9aKa+6wcNvIxDjX51kkaJoDN0nd9cogjg1SP5B4ciRd
gimWNocfJTCTwJdr/Vb3j/An4HFnxi1pCPP7PTf7lvwB9nFXqrwipQN2HGVfOqRNpBlvJJlSVH5o09J6cNfkH3cZLtryYSwCGYii2rnNTTD+KJyTQCn9U1LgmASh3I2S
Mi66RtcaY0yCz7Gxq/dQgZEmvCB6cj+afvRwBWEQQZoJm8zxMW4UKQIE0Yv0qo8gJmlxbsbWxnORFXRSugJcwpreJi5dG/565Q1pwjmXJwbuYyQqVF5M/JfORfFPlZ6R
oAvLtxJG6BvDHMhIWriwmGxLbL2Q0ZFKW0FpFg7/1dS7Q18z3LXWovqQuvMRsYi6qUAcY9nqvzSPPEygbvZIaILIsP8kLA5rrQgFPww10M42e2QiyzVcEmraG/82ruYi
ODxZQRmuUH1fbGZhwayK8lhswVP5cqq5OXW8l5KtwiHCnHi3P5VJvEgzA2A+ESWHgmQdMFf4PIODusGToR57ied8jtRkGiXNoP0nV9EfG5txrFJ9wfWl/sdOC2HjZxrh
MlKO26wPr/hdvMaDKdMGZnZzuXiDsQQez0djfZgxgCOD7tbtlAz0oyO0X1hnxpHL8RO4MPymqrwFvU81rUqGFOCZzQSwj1+dSEBwkQrRqb0SRKb1ckmuVWYo7he2tsyo
BkrsY11ZLrYfuNCi7Wsyp5QHQaYbbvQf1Pt9avxEeOwHF9R+VqtndpOEyXql+XFG/sNfV7e8ea21WC5BDNjozKQZbySZUlR+aNPSenDX5B93GS7a8mEsAhmIotq5zU0w
eadN5t5KlcMptlWKP+NtmzvJwcUK1fmyv1mnIKeM1wMo3MLuRFMiUPlsCsrQyQg8JbmQkugt7hq74NH+AL6kGtWwFM6MEXLiEXCqY50RIkIvcy7j6SfxsM7BElXAQiMH
yi2VO4Ic6LauTMT/37dUxLtgiumYtqBMAm1r/56MFPtJsZslgC2/rxNspTt0Cf/DDbYsu7C9SF70UGqlhG7LBWevpbTnI68Kf5EzrxqL5D+XDe1bhwpE0WHI1rz25raz
rqQPIMZHQqeI1JCudQ4FYqrDZeMV+KFzooYvK3+BMo73PdrOAIGgG4Wgmjqx7s9U0cefRTBG29YgY5uhpzhvalnBZY429/EkJI0DW89m6fa5FS0374ONPs6qx9BWnKWa
J0PJwPUPeLv8y+bGbBqdQqWwCp9WAWYfdzC0qboJSpOXLwVWpmw4DyZwCxq3bnwn1opr7rBw28jEONfnWSRomrx8ELaoeNaS8gD3qvfVltdjfSZrL/E0h0xBch3kOtmX
2CTB9b4nWUj44cpfEF+iAiqnIn1Kq7sJQOxaiJUBKC3yWHuWgqB2+Y+FdENn9epTLUSvHxUrbbkgWUceZLlP+NpWNARtEkeAin9W6yEcSv4rfAM/vTL/TrHJ69UGgnwY
ub0UDZ0qTSOSFWXstqmntO2sVNOF7qDco8Z2GUu4QmnbvocnQUV38JKhbp7/Pq1RmODE9I9RzvZR8FXPZk+VCpoRGBrQvMx5N5cJzccovm23mThM+jaRG1dPb3U7SILi
/9a/QIg5INEkv7Korprnx35wu/Y1vkEbxK1A3sNb6n7N3blL0nymAc4S0qSI7CNbX7aLw9jhUcNJ61wZcmMaWeiFZWJ2t8GVUISjg7vtJ4FwfVqhJvY5PyG15vYNdqJP
ppnBQG1zgRb3sn5BGOU9i+dWdp1AzV1rdoSslZ88oGHuv8wdDMWDsStRJ8uAeuzmJbmQkugt7hq74NH+AL6kGhMF0qjpaNhkbnBk1+7DUZ3CCfOuAIN54jIyzSu+wbTN
tLSDYa9rSXaFi8kvWa9MaOfBkItCV01+2akrzZaau53kFynLkixMGUTCoOu/MdB3QBmcttR5f6b8fMwh9mAEuQJGFYfNUotiKuT9H6jB37ayVPe4pYOEFSd9eK81DIcH
Ns+VYRj0vJjm8rcE4ogFB1Ykwucnl7aE069OEot4gY3bgU/h3wV8q6YoCrDUe0fS8AxPHfjynPXC7Gh6EPS44eeAuK26k25GtDt5PaNaJ2FkgnN/BsKXNAdEb3z0/FKt
PBrGQG4O4+pZFgN9+TsgbiBcjhxA9SppW271OsfNWgJVnaiNqq0D+6Y/Yk4FaLyKFXIN7wfYGl4+DtniLzhJ//tsJi7+Nwr9lRsFayCmrxF6tox6npPn6JB41lj0ozK7
zKw91Zchd9ucxO5mTFxHHamHZIb9NQbNwHyYvNsnmIySToYhYis6KMk0YV+Va65V5z+SAOsbE/3fM5Nh0Y3Ew+NLxanv6NigBnPrtNQsDYaNbrbtyfQD+yrwgUOlre4j
Fjen2/P16sp0Zu5P1B5IHiRtaB+8XeQexGqz8Ygl9ClKR61hDfeGnb3sSXASWlAjbqAFTF8j+CYmimxg2LvL0UtJEcNucnyIRsy4iot4bWoV7Y/flR0oyPDk50hajYaP
V7pzTC7u7ze3gYoxhbK5PeEVeYBtHot7eYFbO3lBiAEoQiFJY+vNcwjmaDCsyiI4dr73VTVHIosB+/uVjfUFqWth/x70N4C3Z77z3It/Ew2z6s4HvoNtgafnSWkCbwbA
+IYA3z0MUUvvQZH1TtrJ7dHQ+sQ29XlfBsFL/Z1DZHGv3SXhzC33RTZGkRYGVvJz9r8QnLJHonaK5IFgw+qI37m+9X7YxiE2qmA+6l31/42T0mwGaq3YllErjRmt84H/
RikVfgelBrRQG3beA4/1faQtlgvq5Hp/YwOX8NE5+nlLSRHDbnJ8iEbMuIqLeG1qFe2P35UdKMjw5OdIWo2Gj7UWcDVdAIwafcAmvCURGcrveBTQW0n9kFpGuuCuZ2WC
ViTC5yeXtoTTr04Si3iBjSBVj3lcBU3m3hELYtC5eM0fnR6LmagJaJ0fzV6CvWi7nRu+6k9KS/9uQT10PQ6gcjnyYQ/qbRXsentXWXZGNFwbUgrDlo3tU/IKmCcKwPbh
2/bKtlshAIdjfLyduhFtRqmHZIb9NQbNwHyYvNsnmIyflYvi6sZevgrPj1IRaMUeYlcMZa+isjrtitvtb6YrZBRohEeLkrWPSRsNwhsVCRYbf+rjSC/tHr8PQDyJ9mvJ
Fjen2/P16sp0Zu5P1B5IHgd0mLnRE8g8cTICs6SAM7j20nZOVHssR9YAAKpxZGDc0lmc7A0nEIGIAduAw2nl9g5vJ960F8pGb5RFw6JLVPbzLJup3x/2Z+xjdyymrXEE
qYdkhv01Bs3AfJi82yeYjC+tCmO1AVIbelFmlJiMDoBu9VEo4Kjh+mJzrq/o5trIy7itz4GOoB05NtpY4sI9I2NTQbkiXRz7EZEB+ZWHhkmDhffmi1rkcCukQeMZ6JAT
K9CzmFe/IxyZV/Qltvwax7SolByl+r8fvNRgshaHl3tSdQDfLooTLA52hoMuKqShViTC5yeXtoTTr04Si3iBjSBVj3lcBU3m3hELYtC5eM1srKS8LD8AxcFcF3fbXV9g
8sSi+DJczPfKbhBpSc/vYnq2jHqek+fokHjWWPSjMruDhffmi1rkcCukQeMZ6JATK9CzmFe/IxyZV/Qltvwax/M5mg23rbRfX0DQThpUxsLjBDAP0v7gb8YMLPMiP4Qu
VZ2ojaqtA/umP2JOBWi8ipI+BSmTVyewGOo8DSQdOzwhtbXHKo5V5OJsC1PoSO0GUXcgbq1/1xjMl9zk28e8rBC57RP9wrCE8NB7U00le2gIaxOmnYZz1DxyzXVloNbu
NqpSj8ue9wBTnXr2BJnmPgFFPY3B76rtIGQEkanXBEGzPNrcS6g3UliuSsyeYVAkODvCuSF+USxIDvKS2uNWzoJ7aU6JMF51pMMAFZ11Ma+xP98U/+1tt0hGbL/QLBQL
qcFz9YAeIlsG+flXiiINJpC9h7GfKGP6hvJhGewQW/PCSFOh3NEe1rY7BHtMl44Q5nHFGX+unjc1ax4939y0IrwqtTlq7yRgUQE/kY33Y3U2z5VhGPS8mObytwTiiAUH
NQmFVZnaGzjsKIWUdvltIHQLnS9sshttx+xnxp771SxY3noTX3DQaFj3JCbakpvdfVswNDWf5n2PZWs8IA2YolAL+Z5cA3nJRPxH8FkO24y0ODvGffJuDJBUZSjzNTmW
HfAiXCTWzr98WoJGQFyE4pKIx+sMNtiX45Rd4B8CGqd/MV4/9H69lrv6Nf4zpC75kkHGvzqGWf7nji3hZ/0F8LosbZ9MalzarQ6lj348B8Cw+c1TIqcjKdfvLhFY3DWb
AFZND7EBl4SmnJSHvllAD2QcArdIL04+dEVve659OAMtB0HUMt8+c7NK82ThujAderaMep6T5+iQeNZY9KMyuz9wCAcv/tjBZRPZO06Kmi/8CvFL9nXrqXZvAioIb0/7
16lAoUCC84ZXuwC9Lq7xlmQR+Y1HwpPIdou2Kpby/MWp18ozZVxFWMUC47VURxVFKQEBXYQKsmGFb1m3KoRcd+Q859dZND6rVzWftf1y8ccRjFWQiGAqAI6N2Z2L67Ld
AcTvF8gwooMKmKArv5m08HKl8ejkEAs/XoQx906LEuNfB9WYCmClWW0m7Yp5Y59y1AfhhCzuPlQFxJgVFmRENKAFjtnM/5OF1nbJ9w7WXLmPD1iocO9zxJVczRPNXA2M
K9CzmFe/IxyZV/QltvwaxwxuUhV9r1RHmFUmgAT32Y0sVA3XG3t1nTnI17lj5RQcueJlKzaIKLtl56xGghAkVJuzlKcqq/ao33z3tuzsegKUB0GmG270H9T7fWr8RHjs
BxfUflarZ3aThMl6pflxRkQ15dgdB77IdQXIx51UHkLLiSckDfCWPE012qkER+dtMgPaj+4Od1vZlefTVY/MEkOiR+9F8EhoOBexeVQbsLtAAmeZuvlGULypS2cLqdso
qAiFsBwMgBtoaRm3YtERU00h0kdqwlyDGBz7jGDya2Y85WQAwz3cq+KebwsDGQdkDyZCRSGpttLkjSn56ka1FgWy6mnX5bLUIQED6TkreKo2ZEzvdtfUcQGIHBJHPNiH
lQIlSVckoGEJdMMz+EwqIsNmaWFzHit4i2RYhVWRn/K5p4nkWaVxLfYW+XY2kBIoeREUKVUcfwzwfvZvLEvl3Fv/++9nDYTaN02o+fBUSd3zIMPXJiKCUqHg+lMni+ek
+0LtBSOo5AEY3c0dEKkl7+e0DZGwhOEAivViXLFX34fFwci7QFNmvMAjqQYI4/4AfdreX92L2lQUEGkisOren+k81wjj8LtBod+tF+N7PNkxYQwWtXhY9pnr15M5PALm
BnA/5HWOjZ1e2+5YVWLNR6vW4SkdenVPJcg4bUvPlBwvBNOBjmTvYuZvwHgFjcnZ+OJPLAwv/qNASAGx3buDiMSV5BFwv06UCd9gAMfvGv+pkmQYSIkk6EkQ1XE7u8ja
NDBlyGxsDpxRh5B8v5ijML0GF3ONIjvhfsHD3vIL+lOBP6NISsTlSSV2qwenXpHU+R5NkO8zZU8ZlOnZKfD5miBUvZeIfI3PJPE2Tgni484Fsupp1+Wy1CEBA+k5K3iq
qildiEE5VXuJBmJGejlG/hcCOsRK2ieUSVNJOsv4C/jDZmlhcx4reItkWIVVkZ/yoyNMKr+pfXDmR1CW835dLPOAA/1sjmB5Eq6lT6E4SzJb//vvZw2E2jdNqPnwVEnd
v+yCEO9TkuHVgBlXqh7WF5JvLUKqtLcymscnZT1r+ORb//vvZw2E2jdNqPnwVEndTVYswwCCNDf0riUXmqSQDqpbfpzduRcHlTFrfL0GRu1uKwaDh3ZQ3noyc9szit1s
4yoozviCjXGeLMZUWqyjd63MInXKMa/OggO7bv6XjFaLoYonKASdP0EGqVwcl5mL5TjcjXTDoqUfyiNdncF+w+vfcoqfSa3tjQLnYNAEKqeH5HGW8rz5/+wbl1Btqy2S
hxGCiu9+5I/tqHW6Sy3k20g3ZTPo/GDb6GC2Tm7XjWyn7iQGf8ebPMpwOzk2G6triIIY9lWHyAFGTQvwncfOp3PmwdHnOEQXlKBKutzWRH304vs0U77cmzBaOEXxhXEf
9lZDInbDnN2z1Bi3NvPgygdv29sYtUuRoFLc2Tp7ccAe9MOOEa/X/Hb/Y5V4Z9GDB5yDm1PA0TbM2b/4kNuYdgqxhGQLmxt6C55HYo4ozkiRCNq5/BFBwevjBelJ3qrk
rBzQatRW9rPm8Sw1zfJs3/hBNAzusx/epL3pXmlW/zqV4eD4M93UTxsFlU9U479fxGgymJnTHATawg5s/ZL2uAcyf81pjDhLIQfJol2LGjv/tiTBoP/iygBWN/89Khlq
LMXxpYHu9XgqiggKgkSr8aKbDOSpyzKgvP2NATmVb6/Ya0LT4tetXzeuqvfGNQQTDBM0oVPajse3bjTzYmfrp11/ZrJm48SYUmL5l++echQ0aG2PswtQyg+YBdktcZIx
KQgjtmkTmNdbhmVohurBUBCRN99GS/MqArF36CxjeQ2kiaOBvYsf6S0PrQctGrNxHJb+VT9VR6bS/DUl9pcT5woXN6LI59HWh4aJMK590agLs0pB/FeysrAMQ5yqG+35
gZC0IG56Lcj3BVGkAPWLisqoWgMX4FJJUiLGANLwMt/zLJup3x/2Z+xjdyymrXEEXnP9v76gso2qYPiItTeJ5RzFyrk78+15HLA2MVNTjHjb9sq2WyEAh2N8vJ26EW1G
lHO1irF70vjlvf9cC293HEI2EEiJpuKXBc2/UVAfYEt+DyO5Ewb9aJ3qo59ewBzneraMep6T5+iQeNZY9KMyu8G4Wh0ujd7GUdpLSEQt/hD8CvFL9nXrqXZvAioIb0/7
16lAoUCC84ZXuwC9Lq7xlvXq6gVC8SiRhvcEGURd9XNASZuslT5hhBN67jA6A/j2pC2WC+rken9jA5fw0Tn6edHLTDNb7oBH6UuUodoeaGfb9sq2WyEAh2N8vJ26EW1G
lHO1irF70vjlvf9cC293HEI2EEiJpuKXBc2/UVAfYEsjZVqYCS/QIME0EkbF8HB51AfhhCzuPlQFxJgVFmREND6AJT6QzmTgKORQek1/qsikLZYL6uR6f2MDl/DROfp5
BSxEeZmS3NL/BKw2+tLPRz+r9esPW31QZRJSvwlbT0nK5IRA0pCtUUsOC8LTE1z4gKVl5xXZdSn+nQLn5k9YAyl3cte2DrMEpj7DTxSB4OWUBU+LD25lTotcLq1hKrXc
LzbURULGr8OcGsHtJ4RPZz5B1hlcM0i2X4Qr4iRMCT2UQakWoxTwHXjA1UVKJvNPHmLr/qDxX9jNe9NQyZ+EhrGVylnVnlONkmP6VF3gos9ftovD2OFRw0nrXBlyYxpZ
WH2W3bQykNN2RhhZBTXN1DY221F551d1nLF/lIuYe+AmvKmssOx9a+N30g5oyxGok3Agi0yDRvKGHNPfMg/tlAsnmHdx0iEYpcAkLfUfAUMDLqaTsAHpQlphxclpFETR
ub0UDZ0qTSOSFWXstqmntNndShPzkLodk5RZ/lGYTtQ5/xkO1Fhr5qBMRXdfGK1/yuSEQNKQrVFLDgvC0xNc+IClZecV2XUp/p0C5+ZPWAMblwIAs4wND5yKxP/GrFeN
cwL8VlfNcpWwgDmeptDFu+6v3HwSFmTpGkyILUF6Ue9ftovD2OFRw0nrXBlyYxpZIZZ5sZSV9+dff5XDGsz/dgm/j9OSVTQIJrywRmcpuVqpR7xlhUDHNcxE/op+sFGL
9+Prl8oCYHicI4s1G/PzMj+r9esPW31QZRJSvwlbT0nK5IRA0pCtUUsOC8LTE1z4u7vx6ForocW1eYJIKYZHnRw9Qim/2EGHqKx5KAPymwj2d22BCzSZkAkBGWlH5aTE
cgfnnStw2Qa8FgmCYKnmMdsA/fv2TCb0eNywn0hzXkwq/6crEUXICvp6htTgGVJn861XpeYFOgLNe9sb8Dv9TJB8q23r3oCFV+/E7ceolENftovD2OFRw0nrXBlyYxpZ
IZZ5sZSV9+dff5XDGsz/duJ3yzj6WxZqW/SaF1aS6b65vRQNnSpNI5IVZey2qae0WhdxaNCiCa8Cgaynhi78Xy2eKiBZE4tYPKrst7VjyC8Ntiy7sL1IXvRQaqWEbssF
D/kEkXYORgkx9NcYxk+d0TY221F551d1nLF/lIuYe+DLiSckDfCWPE012qkER+dtk3Agi0yDRvKGHNPfMg/tlE6Hcr3pkc0t3s9NlcFHPM73PdrOAIGgG4Wgmjqx7s9U
1IIczQJjrDJNozHl6k9WP78HW2ZxG28ZsyGVM7fqKGGG/nAtueWTRmVxh/d6i4NsKv+nKxFFyAr6eobU4BlSZxN0xlcj3UOp+29RoO7862s84TRRo0qgqDbSzqP3QANZ
X7aLw9jhUcNJ61wZcmMaWSGWebGUlffnX3+VwxrM/3YJv4/TklU0CCa8sEZnKblaqUe8ZYVAxzXMRP6KfrBRixISu3/ztEuu6gxtedyyb5PLiSckDfCWPE012qkER+dt
mUadK7LXopjkIY093aFmPw4ICygt3vygLi0PDqtRoygz7OSopDMWJMMn4ZSMK14bmrfMFIFeM9TzU7EGCvxfJBaW+ksxA2praOjnY4RtFNpftovD2OFRw0nrXBlyYxpZ
tQO/tHugf0n6HvmgSY7mAZwHq9O1TKvpBANWVIO9bA7WimvusHDbyMQ41+dZJGiatBstzJCrNN05VbqUUq/97XeMGLkMat7It9uudHH3jNfsTHTqT8CcSTqTnCxhfkJ4
ByGy1sVuGbC5FJJFSouDuPn1XbxOGQ7hTjMgOs5xF/8anH/eVO8JItCFLRknIwfiz641gvotR3FK3rfPAt6ys5LBeB1a6ThdMgjZJQsVP7tcZXtgRQ1SqqG2s3ELcd1h
sh0LiQyWxY0M7jFTO0ftQ/tVRPRspbGH3ATepu0KOsgltb9q1QwfPkDWNkYjByIVlTBIreUT7FmPbOpfcIGaXQGIPpP0NFZHqmvV/BD6v5v/LMtglCMaTBxHrAt76svp
GEkMWFMcEpw2+V1EcJS0C3N0Rju2zlUrHMLX6xL6jdRhbCAhlnlXMSGon+jVzPYWAw7ljPmZgskBbzOLUb7JlerZ7QMfrosHJWLfJ/VBa2cSYew85/y4z8ERXbmivYEJ
v+jc67Y3nWr7tAbGyoWT7rVTjFFh1Mp/fS5J456Trir7VUT0bKWxh9wE3qbtCjrIXLhJc5AGToE6E/vz5jzltpTIxe7sUCkcNxl6Xq8h5GZXshmw4x3PZczcUKbCrxHq
Q0YBvFhsmIqjWF64RIJfO7z0VgeFBFriJeJG8vOSn58hRIkf/Asfvc5rtzR7gTI+uFiO9FbqWdsqf3ymC89kDmkxYyYC4/Q1NP6qexaTzlH4wgfcPZIgSJSLexOSJNSb
ieiBCPjF0O0RI49RX8BQj9SjUXr10M9kKfiSFBu5O0Rd7ai9VclZ5kSjF7cIfiaUFjIaOUP0mH1+27aTPlBSculMTB+cSskaAf63afn1FETQo7BL7dpN+OvXXz6L/iL6
T51ePqpRpqltCE69Wav6kQQbVymYzefzTCJYB7wMLVsx36/Px6mG4dRUY2z/In12Oi5tpMU10IHGNmS436I3cvCmyanZwheTCKw3v2ClBGckiFFgZ88TlzNBXnPYXASg
Az//jdMWyssDUi1IK6hj2mOsqWnpyXlEdh5xOg0Qv3qqs6LkGqhWxIHNe7oDoLHUex4HpGEKwnHZdzzgXglhvrNVx75SO/dP0z3Jvx1y+FhX507Di/1b3pvrLNJsLIaO
koE/FJ2WFQKPMgQ53+GkxKa3O/PbpCqNcO2h/+xiEQe/0DYYsAU+zkwlIAorbb1xV7itL4nAHCp/aTdZBcgHk6a0rrF/bLEG8zmInajKnb799g62vJrpJ4+5F2YZNsqZ
bzWnv84gcdOoKbsRoRBMflCZ5uryw8iKbKK0t/07Kwf0M5hyVzcqCDpmYtF1nNWUx7SR7VLdLg5NONuDvCfR8XmDVesFrY0WeZGaiLEUMinn0JI34k8fBewW9NG6qz0S
xuDRhCoZF1D2iVyLPKCdT4IkFMPDC5pSwhzipB7HMwO/ekfy6LSld+shoG/iPJTQbvVRKOCo4fpic66v6ObayKSt/CqdNisoWccltHEtij0uzClQFaq2byp4g/CwVaZD
KtIWoBgGb4FPymKFHDodCZtgACEZ/iWCwdQBQWY5bIzV724Tt3u1C6bR6uvXwXDT97ktI1yD5Psmj3c1Qp23aMC/2P5yyD7PEakQ8tbcaQZ5HzDAD6H9FQI6W7mAbm6F
TsYq4pFdjUN2wimFCUbWtBobRhkVlcqDo87MUSIG5PKQjPfNQlmhJVU6NSkEVv5tHWeA2vpjsn+7itvFWz1xWeb3gw8LuFe2W5Meo+1ql3vcQwtgh1dHgmmYMGaYnYfZ
6GtxbvwG+PrdQAPXKbRlHa5xB8MGyTUz0Tg4aVH9rzITW1GnmbpeCEjd/tzqM/nI8nb+gZ9io6VhcZYgC9AESUkIvZgjFNVGshXb42dfLO2YvA2DTnUznMe5z3oUcl6c
4uy81g3am4KNGpAqxlkPxw69sdyDBv6jSse6EAOlo1VycPFY9ogtOHx8z/sVKJvpo27qCgv4TIhRF/NawqePdIfP9sgs5kX5qyLWeG4KrOYMtcPzchDXVke2ap1T652S
bna6qC8C/fvxHNNWE0FCjYmZg5gT90Pksa9Y94TzcpioeL1X1FNtHIwNIA+phu02ubWK/zIY4q5hNA/u9UXlWzToUpw6G54nDu9PBn3naGX60TD6ixAuQoAnGyoyvt0Z
8887u5JVeLia+DBy/B1vLLwYNMbj9ezqX1PFln20MxOw27DseU4sD37CTI6D63v53wS34NhpZFYDo25QK6Op18cpcxghWcg/rh5aW1geknPf4bTE4foL3uaXTuVymKIW
yPkkRqku6AypZfR+gS24+tbc7DTP3Zb1xO+MxGVGUcfthfNmK4soGVZsYP8ws71tRFhsL+xKoj4H4xv6xH38oe4yD51jT8BWlwKUUrxIiNaYaRMyMkJ8oCQ+qFOTVPDl
xk2YYG93GLFmXhCUaeRE7rfXCIv2ku9q6ca7wAFnxGC3qVTOGAGU0aI4L4Z0jekWRnbv2attIpjNpKd49EGO6eYuA0N0o8qI9ZbccPZIxT4pOGY1JRzINgOl1vbw8hzw
vRe/tWseFfKxUqC/op2oSDXOyIt1O64NNU4xG8+V1iH3rUqOOiTSIdhTIMg5HVium1ckvSYxOoJFvKdlLlFDlCmO/G8ONsRIAQfXY3ibsLYGKLH3IJQ3Dhg7bCuBDGKM
peupHKjY0SuMTsjc0TQLV8UPesi6j8abZDsa54cs8DESetL08PX/90cT/SsxT2S4bDnXjMPiOdR65htcTFryqPKdhQTe0sz1UxiGLzU/u2aIbo6Mhah8FCquoiMKRB+y
3pAg7n5f0XjuHj73y5XghNn9uFmWU4jkIOfkY0OppemchnLUwPJA9Fzm+fkQqImIdqGOxyAy6So8K5gfrHulpI6fx+HMXh5KOiTKtRl69lXw3Vo/GZ6/DKZ0NKV/Ae9Q
/VIsN7woryrYOvMm7yHvKRTgXYnZ7QvsWoAEzAnJvdP5/rf3IsZMuKCcZsfoCDzfWKIz9Q9vwx4R442Tc3bJr/MITLWjG6OhHQpfcwJlK1IUFp7NKU2I+DlAE+pzJ5yF
CKqwsWoTWZbfeIjLPTsOVdCV6AyJU3lbjIyO/1jF7+V/MV4/9H69lrv6Nf4zpC75IMCJDyp89Ap4MKvdJT0tIEuxPoqnq4LRhBIzktBIPqYv6zNRuWrjZDG0TG0Csfu5
vSf/byC2P+ycXnRtYAbaZliiM/UPb8MeEeONk3N2ya/zCEy1oxujoR0KX3MCZStSXElCRe9uXs2HyW9fk2RleKQtlgvq5Hp/YwOX8NE5+nkjFfpq6BOHnuVKGOjxEY+a
Ns+VYRj0vJjm8rcE4ogFB0PaYZn+AnPy4xrt2vPc8bf2tuCZV1stHEopAUgUTyicoAvLtxJG6BvDHMhIWriwmGxLbL2Q0ZFKW0FpFg7/1dS03LE2wOx1NnX8vG3wDz9W
Ym7g4njev+mCxidod3fMkqr1MG9bNrQmD+ryUSecVUoeZwTMC0/rBJXC5QKs6vNwf5jFCcYJ1wAnbhaNbQXBBCMlg0gQek+Ye4pKSPMNXLSzRYGji5dKJIsIC4XZYY2B
m7OUpyqr9qjffPe27Ox6AkWrfu8kUs+iUUqKsOsloOm20xbNGIzJP/sRi3nPdyxWLFPha/iotgN3CqKBzg+Bwi/rM1G5auNkMbRMbQKx+7m9J/9vILY/7JxedG1gBtpm
WKIz9Q9vwx4R442Tc3bJrzPuLpGONsTGd9cNqV3ZXO9LEnQNTgelU26eOw7MyC5/4BXXffItfpenlpC7GzKbaJAMgzXXzJ9bzotSH7WNs/qpc8cXF8PKZWW+LkYECC20
GkW/oP87STkoPtvsGDAditpWNARtEkeAin9W6yEcSv4jEDDPrF8BbmkYp6N3L4hO6OfuNeETtnO/tx7QWTsvACEH1QPgeVfctdhF63fW4Ls/A4ZTu1W3clHCz3yD/Nyu
Q9mbZex0BDPjF/m5QNG0QFuZJzrw5l6lHWUIoTD3aPmHmCcztPNykKPxxY8Tv/6S32Xelm71i1zWqiCg793Cpuvc+E2KCe72bWwgDGu5QtTIq9KlH/WivPmt5m/Sa8Sf
O3ST8jTIRhS/7ybxtPk/Uxku4wzLqEALDn3Yz9yPsLA/K7jXy2SI1BxOeWBKi5Z7wlAWWOhFEZIiga0Onzcbc26SmQCPjN67faQ+Z7+3pEv/J6mDU25XqLk96UW2DosG
IQfVA+B5V9y12EXrd9bgu4q7j9yK/UP2aT5s5cKJTUnZKSsmDjsFK6tA1+rHzueSIQfVA+B5V9y12EXrd9bguxlx5I51loo6280cPE1mcPaTtSLnRRVzXi3B4pMkerTg
IQfVA+B5V9y12EXrd9bgu0PeqTpQ7Yr4qc5GM7izuFPDZ5xQL5kKHeOshWZq5+dRIQfVA+B5V9y12EXrd9bgu4OphNus5isJ03o+50EfbKktIaiYgNP5hahY6dIN+oOm
IQfVA+B5V9y12EXrd9bgu53sVE+fhn16TFjDAdIO5GEHNoLY6kPSOjWeN8vPv2q4vVy9sWVIUOX7JIds9QQqTyuveVkNq264gwyxA0I8rjDvKjuxH4PJtzYby06zUMSN
hcJ1q5d9kmKUGKmAw7SQ7vCMo8VtQBySd2OuSvppIZN0+ITXuJMprbnWGD9W4Oa1mbaUhvBzi3Am7waKq+MklcHG2iyjZHQuKlHHA0FtYzwI2CjtFfMxlK9GZ2YfoTAE
ZmuPyHa9qYqctQy9RFYkuG8D/EUxKxrhWclHbt7Pp/4RAjeSE2VMdPXa0htlcggRf1MJAPY6x1c5oaO1N7TND1u6/2kzFHVb4hnsHvC2IjkjqtqgZ7eJ+6cBs3hJ6SRA
NplzELC7jjxrUTmugbCYc643bIvunGZy0enOuwdP1xmq6Hv+SzR7f9AzTV2CrDSnBC0hgrjSjHw0KGxqyVlNs53YnhP19JuUue2sWKfGRFH+DEzpcDxKuWD8bMS1/vZ6
KJZAmmXNqsXbjOtpomcODH9TCQD2OsdXOaGjtTe0zQ/UubFCqeA8tIO4brAr5FW5ZmuPyHa9qYqctQy9RFYkuPclJfdJ3oJmxIBrvpWqpbc3tUitEJffpUY3eS9FJJ0i
sRl1g8bgl5HEBOdtqxaPHfDHiKKmjT0bKw03H+Y3ZmZ1Sb0eT/QBmfIFCZRnyIQn4LO5C3j6oDMHD3VyNeJxpU5Kq1efaKB+LWdllNkUQqyd2J4T9fSblLntrFinxkRR
uWX5oWcf5KOUD247kfe7FLse6o3vzhoJTnDfQlFMaoLcnCykz9dRsMMnv16BP1ajSDdlM+j8YNvoYLZObteNbIUKcBk9ARRHq13dfaW04dDaLX0uxOCoG0CQ39fnSqQA
otWERehLjnODubns+SJzdV/EPZBLsSaFqRyddkA7EIfFwC4WVhyZbaAM8Czw04NxpC2WC+rken9jA5fw0Tn6efeX9mZTVH4RJEKx+/iNkdlfxD2QS7EmhakcnXZAOxCH
ZOzTbdg8qkgINhL8FA60GiT3myxFel184KIGv12c3/k8pcwu1dfLoMykcbZoZd3Ls+rOB76DbYGn50lpAm8GwICWi+x6ZuYlSkRB0ZTmVGlsS2y9kNGRSltBaRYO/9XU
mRXTcmwLEzESIAXqtFoP35PJWoyh2xH7y31BhjaNkCxp3K9W0fgDWPuf0YMo2uI5U3/KnioULKb0QGIp+vLt/8UKWAJ3licKSIUktSlhfbiD7tbtlAz0oyO0X1hnxpHL
8RO4MPymqrwFvU81rUqGFM3bNu0gJLss+nJjcYhLwle+h0oRGnuF/ekR3voYBU3rFGiER4uStY9JGw3CGxUJFnXnjWORigBtaoqglAmZfegwzTrMCwPa0nUafh2QBLA2
Kfd6DfWl2VY9UCqM3eo5GUbI+dLaUrSxUz67vBGeDDVSn5ReU2lyC+Z9nFqq/FwxwEQ8xs/aOSUHhKLw6znhSr//XpYkUddBX+PH9GH6O/hJ1rMB4NHabVxkt1Ud2DHI
17kgvubk5IW1i8AJb4pR/2NrDzgUBgW1GklQmNGllDY56ew9Ur35nBbQDuSE0oWXXX0P5NXEhCbZSs0AJrU4GmrcZp93qo8nb/zHxinHASJCYKF21l5okY41JewekPn1
temYsCWMIXIUmcRt5t7bMyn3eg31pdlWPVAqjN3qORnScjsCnImkkgFwOD3w2PDq5fR8Ah8l15eluZJINzb9ekGLK5xTbco+urrHzHxBfMLE/5fMLfGXQYWTCSuHmyha
UnVg5+xeeQzDhnEoZzhu1IQfP09BZT/4JtSlDQS1nsbSMRig2FWdq9miMjZgoyqu/HiX1tghYco5hY/4wpRsBpZgiTjUJI7Y3AGWPmTw9D12fIcBKp0U6S37ZxXXSAUX
Q+w01OJJfKh1N5LQB6682EaF3zDBZYzFSEW+at6vvielDlOaMNiWXhjv7dgjm4A7mF5lDNoAwOyZc8li3b1ogwlJOvVAx4DtYG3jMOljXAey655qBf1+9RBAOu2vc79J
VAk36FuA/b2Ye1t16DE6ctDzTqPqb8D1wRtgUmhLc4zkI9550O4J5BBN6e4ma/ceS5y0iKLOiisI2yN10KWzlWhr7rN+kiU6cCZFf62fXiooTv9hKAZXc6mCrCuFq3xa
x6HZgAaNkuUZVR4vZsZ2t6p4Ns8TWHOO20kpgxiTjsPQJU+ZqMPNvFYiIELsuzDJLAjR55ZAAvaUG7k8OutwVoFevnWl5FDpSPrPRno36mF0QlGOnp4r28DrPe/SVJ2+
PBA7RfUx3zPNF+w48A2Gq0gXwwY+NvP6S0agBE84fOYmKgmD0V/fG2YsSvsVhn7QHs6yR2MreyEtl9W+DKfvFwy0WMmfOEX0fUJt0LQpyftNadQMMePo7ioUDoFyNAky
juIrKsTnJIIcRh7idmUt4bBNNf84P66OQtIWTuFrEDN/+ei9tTf5f9DOQlNhsXj/suueagX9fvUQQDrtr3O/SetlKtuJI9Adjo0EzhUAi1ZBA/po91ZtDM0BC+BrNs/d
v3t+q/ZX95lLyrrOwLYnTcR45vQpgY4s6RRXsXa1jnYLga+Kz7aXrouCdw+jDBowkJCTdROZ0SLlAmOTa4bXH+vCizv6zsjAo6SiHxbyXLjuNuLte4sQVY4/hXjNiGqa
kF2vvKjpSw2gVf1QoPTmOuoc8uNdI9ejxB14LTCCaU2VudZglfS0dFeSQ5L/crMDbDhi9KpRVT+7MVChfM4M1q95XEvJ7zGb4uiYS6UTjIIBBRV2Ws+Bo4nHMZSBS5mo
49trqAwV4HgxC+eaPU0+sPz0yyP+lSRUUN/NRY+DdC/uNuLte4sQVY4/hXjNiGqaXB77y+RuFwYvWxOJr0XrneeTaSSIlTTW8SqbDQLXv7P9e+jnQzTUiUeflyUE4Iru
gwhurQiqtt+96BR1/3/b0xnYz8TOmbJeSUIb54C9YWiaxVZ+5SHsfw7UQtv1LQykMkYpK0i3Voj7upHo4DLyTlXqMo4NJY+x5m510pRtExDjBP7wYEJqV5SwNGtOcT5M
vHzMe/bZXpDHm0t5q7/yvXRCUY6enivbwOs979JUnb4XbguPVB6eOyl4ULEV/mpRRUZ6gzhuESLeKApzhRGi0hytFCFX4azbU979f6j70bXIvpPvM81OID6gLx01G7lc
twD9/NX5ZzlxLQER/aVjMKmsxJn6X3C0zp+pNRsNHGATBCHC3aSIo7UVR8LnpZulUPCwJC29HD2RIYD0N0zsYRNoG5EqfXDlg6uX60NoJmR+dfwrM65Pl9ZY3v6PWUlQ
YpgBPjhO9v5c55v1TFXM8lwe+8vkbhcGL1sTia9F652uhsV+kX+i0frmKZp1Jj30sPyL/0jXzKj400b1Q6zd4PeQ0CjVHslHmf3v+5SLAD+Vj2IDOQxi/KCJw/fCiCGM
F5VOhE40K5ZnGsKz78fiyVHateR0MlYihfYyuYpXcoyQJfuz9l25zJSGoXD3EyDaILVu0B6+OWAZkDAJIFQ+7XhHxS4lNp6LPf8ACmNA0LA1hIWTrM4u/0hBmpGCEKaL
m2wIoewQttL6sZ7PPKcAM/Msm6nfH/Zn7GN3LKatcQRH4BwiGjhbw7o/UHkHiY/cFipUp+uVqBKEx1gq4cmyLlBt/c9H4XmOGch+RKCKjwL0Z7GNCIlU2Eyx64s/0Bdo
4Od995wvSE6lECLe99i1m6SSDGIdx0i14eTGJhgR0o4p/wHOnMM9JEDwFcDJiC2P6jRnUWig0wvyzWx5ZMMQ9sBodOORMwBSquG6rjWXdnUzm3ztpL50qsvTs/rDWVTS
akpi9IRrweaR6wckoeXAaWL1YuIbEmM6fietUq1GxGALiVqO8kgP2EOR2l6i5aGgKGzcpjEIud/pqyxevEQ3MT7j3hP6HhR2SsNgzy1wpbQ5N/7C0OLq9kI7jtLiLE1y
sbQImGCuFPwCToQMfomL9mkZ6qJqSe+oLwN+jzjiugBFntxJ7H//jUqFIHzjlm0K7TxUbmw57hFNicgdD+N/WMeDmH7lgKHdzf3dsp29G9+RJ99smvyL5akT9B8FYzE/
u0jCBdR9OcvpyC3O54HixXH408oDHgZ2uQdpd4cr5A8XOUb1yOK3v7iCNT/08GTxG+hWw31PRiCFHfcko3CwnBUnoeVfhBVwulA6AOXfje0COjaZ2TbtyVl//sKlwNMN
a0wme93LtJhT0lZDSJ4KEusLLElW8TLOJ+n0cwm0qXfXoZRGbw7ATog5RtvNpjMte8VKOYOfFyslu9gZq8zppu08VG5sOe4RTYnIHQ/jf1hnZ9uN327Wjv6L/9QKFmJe
udC5HEbcCSpevzhbRtxG/fbdIQva0BXfmYlBez1ArHbc4PJMLifBRX85X/2tlJiZHmRvljuu36NbTiS1CQuVtNcXiy0f/e8+iUaeW5pk2h+hdDABEO/71Zr53CwSJ0cZ
Gh2iN6hazAXHcNs9d/e7JlaJe0oe9/TaOHb9ivJZ7z5YiMhRTUmQ8pJs3UODS5PqUORewbo3on+Xhzo0whTZWb0LGRXFa3BW3VqSv7uiJRQXOUb1yOK3v7iCNT/08GTx
ocequomyJbI+kWfL5tcZCIeuIqBXf9VBHIsHcTDX6lLskZKwSb5o06lowmwb8ic2G80M3D5xivdK0h/9qK21rOsLLElW8TLOJ+n0cwm0qXdd8EG7COiiZnZfxpwejyoW
MgC2WV3HddUbguAL4p/CIO08VG5sOe4RTYnIHQ/jf1jM4PeJh7oIMfuEZDi4G44TZqfSTzKMR43PwB9gjX03LndbhWQjVP8FF2RP2hHHWWwsu3I8oTVoIseaSMhatMAf
HmRvljuu36NbTiS1CQuVtJ5p4dPECIQoQa//oyqpWmP/C1r9/UQsp66JSqHfbIFggUaczVbO5npMXrkudt9MZ8vLmpy+l/thlguhtPzxvODrCyxJVvEyzifp9HMJtKl3
4yRFQpGFz0LG0djA4Fj5veOeHXDvVjh0xNDcnU8vlbh6vPop35e5BT5KnVQLLf6Txr1XNyJJpCqfSH2/UwR71liIyFFNSZDykmzdQ4NLk+p9Edjd1oa5x7WJlL4D8KCn
hfOpekG9rasg6a0NyWiQFRYqVKfrlagShMdYKuHJsi56zf/aKHZAqrXNhIm/YlsqNorU67fgDCOhZltNLSfw8Af4gY5+rkNx/0aJhHuFujFkL0Tkbq7tZKEZftQgUYpQ
Kf8BzpzDPSRA8BXAyYgtj3yT0VCEZpdQVxYDOOjIMe+WzaArag9nvtDeWE9+FuxpuLS/juvIPIW5iN0u4OQedQm+2qKb996PhaSmctQs2HFi9WLiGxJjOn4nrVKtRsRg
FZFx+y9/E2bPrhfcWY6On6QFGN8t8yCxWuQK9acbzbR7gqwTs+GGwZ2ajlXjKwiZddJ6LE+qXLPJLU2otAGn2gcH6ORD3+T8nqgi4Idg91uk0dmcP8WpvVKhPdYnBSO7
jgvPAAWX/VM0ZZ2lG3R1F8XTavLQIltphKVE6GDEgFxys+xIxtJg6c/l7FJlQPw2fzFeP/R+vZa7+jX+M6Qu+bblQnBlt9pAJQLoTtd5sTuxERAXZMxajre7wScrDw3r
uvIbpwZXMOGVK/ZveALVitCV6AyJU3lbjIyO/1jF7+V4DPKYEynrTjZ1ltyVPtEUtuVCcGW32kAlAuhO13mxO7EREBdkzFqOt7vBJysPDeu68hunBlcw4ZUr9m94AtWK
U7STCO4qa2vS9NtKbzQrIMBxQBNES/U0OWbKWhwjZAembEJXOoTDslfKYuVA0J5UzwOQKQOJNffijmnep0AUVA42yQU3+Jnl0JzSW6A2+6R1BIt6OZ2/Nc3aBxtP+J49
WhEjQH6uHJE/SMpfZtSqmKQ4MzIv9e7fNFzEV65MEozuApje79qhQ4yK/PE4jtv/95f2ZlNUfhEkQrH7+I2R2UZ279mrbSKYzaSnePRBjukoCQtbeKexfqVWZO2j5LKv
EB0KVN0y1LfptTGmu+Jy5KQtlgvq5Hp/YwOX8NE5+nm3qVTOGAGU0aI4L4Z0jekWRnbv2attIpjNpKd49EGO6SgJC1t4p7F+pVZk7aPksq8eTMRYS+TtuIGmoWH92wUV
pC2WC+rken9jA5fw0Tn6edHLTDNb7oBH6UuUodoeaGfb9sq2WyEAh2N8vJ26EW1GQPwZ2rzsRrtyOFpzXP3j43fe8O6nR49q6ux5wYLMn5DMtdynicCyGzqFl0ujZqE9
NYC6l/FgUt8Zc0TKd8BA9rpjheiyhpGReL0fkL8nq4S5f7UKOJY7Fyahu8HfgIWTbaNU7/3ZR8UZ/oSewGGcyEHIAHhvWFtEmDGf0l1cyuukBRjfLfMgsVrkCvWnG820
eTGYDySsAHA69g3nT3f3agcH6ORD3+T8nqgi4Idg91sf+L+taUCqAmslFxR2ginryHkQF5wiUMozy6tdyZH1gpVZkS2EyyluplhpozlKr1y2fgubrYVgULEIwsMZdDHM
ON+osqar/o6ruNPlhhBWh1VvAUtMGfMejlTDu49G3yjlGbHQ08sbhjD4GE5F1XYQxqffbyFXbxV1EYW+fXLsRZRdrf7MuqoUgfKBd8ST6jS/aMOlIF3aP1r71g64BHFr
lrtQRFvV8gOVev8Uo+ihaV1mMK/yTlUrl4+pDvq94tGxERAXZMxajre7wScrDw3rBdlzFXUtQdBAem4lzNCosVBVDRz30IBa+/yqNQTE+UAHB+jkQ9/k/J6oIuCHYPdb
ZqoZdx2zo5jt9MZwkcpa/aQFGN8t8yCxWuQK9acbzbQ2WaVWZVj0R7niPwEqwNARbaNU7/3ZR8UZ/oSewGGcyJweadVYXnj7kvS5dNLK4OMcJbqe/1Mzpygild/LoVoZ
hcQsWn7x7ufvbz2UZCN2yRAV6EomSlbi+/i4Aqn0zERHm+DTVtSs0ZkCVY8Nh/a7xLWzVDh6Bq01bkn3qblOwGhaHiWR3jryppKTGTOCxqOdDL1PEPUyaHMT86WwdbDJ
rKfAKgyMKoELnYZ8QzQNYmQURRskMm1nvTFOYLTK/Crg7wrXxVfCPACGBhxmS4a7uqgxTK6WyKAbkgC388hoyUPsNNTiSXyodTeS0AeuvNgM4HBNx4vy9tEgP2TS0jXk
BtBUGSlYWlliw6NSTGqssqQ5AzR7y7jdz9u17lMoAXk4S9dnU7k9XwWZnsKggH7lvq3Dm/b51FJ8d2ijZiRXCWzEN8qsJKzGJIsB6xPfyZSW+ccF8F+I/ICJ8UX8WV2B
bNCAdvpFMR6I5dOZSpmpi43faZNa/FbLrY1C806ShYqLV1xfUF04lsUOI3YceuyReraMep6T5+iQeNZY9KMyu9DEj869zF5rMBOp/Y5qptPzLJup3x/2Z+xjdyymrXEE
rV8NP6XakXjvxPYCjOtHb3BMT9t4TLy0CgQyQsFjBDsytMVBfOtexDcXsOGIo2XRfg55uNsFC02HqlvxlLZF9yn/FIfUPfdjBcn/wS4a94ceOKhkH2mT/H8L05IBcNEC
cw1LOSUHjYs7CEjF/nWZl4J5TTLIHpn3eoBQugS2QNWfD9tgbslF6DfKrWe+WuaQbNCAdvpFMR6I5dOZSpmpi43faZNa/FbLrY1C806ShYo0Ljp69eYK+E8AFLQ2tjuc
XkCE/MxIiUru6Xv31eWduTWlq2qrwaRzT/BZ1CY16CAwcMpU6vYanNPACE7n2WtGAHQ7w1ZtYXFOKA6Ekt7mX+FrcpCqdPYIjfBjw+EkxbFu1jAZxkCfzy26m9XA0QNp
ZjM+X67Ftx5xYFavVESedfxU+9y5r1VTaLnM9gqKLrEq7epBC0mLlOOT+TeLRaleyVuFZOD+jo9RXQjaS5pIQzr2P8v6O65JVeM93RP0qAun9lgP2E4K7lhUJiFcuzcB
qAiFsBwMgBtoaRm3YtERU7uiqrhQb02P8bhWgbgRClAFMnhqeNHCb39Aw35VvwCzh72HGo2jSu47TUz1v0f/zobfFLq/ZorJu+Hoshm/r5foiyhqrXqj4lmGkzJNG1C6
oPGj9Rrf2hmwkJ7mAkqijbXSm4vqHFF4U8FVR5lR4CYw1k2lMgL1/lHbTvsrlvyze6uYEDGBCeB6jVOmJepGO/iQaZ+P4naHV64HGiCC37h0VxGRyDWVPFwZZQp0C3Yz
2M6IhAAwEgmX3oueJ4tLoKtboLnBbeSEVn3qfWnBXIjHaNQzaKjLfSkGkxuRzrJiZtuwFZ+FiwErjnDz4XknxlTR4v5Ep6FUBegcAlSN6DLha3KQqnT2CI3wY8PhJMWx
ILn6QdFx/3namTzE9Rr+9k+uTFdqbWfPE3VgKOG+5lt5kuGBPqMBzvcw2WJkFXOA6xWoRdRC/LlZRpnHwvz3bpXgx2KhgWlYfuGQK/2ig+eLXVZHhtiT+/pBCzv3nfXC
YjKsYwkN5zAu9D1zmaMU1M9f4Q6BwvXVLDL406NI15Mz/P9/eHmim/9eFv0YVtu8BTJ4anjRwm9/QMN+Vb8As0Xb/P+AhdkpXJGWjHg1MmEQWOlLIAXE9nd5RltGL4uA
EMlLTKuBjfKpqAjjeaw2ywg7ORuWugRIbXmXer7Z7REesxzhd1EzkL+7UPQKI2nbZBRFGyQybWe9MU5gtMr8KuheRmapnF2z7PfGZPTLBVnVttqOoPusgSPNdFHpwRf7
K+xCUW8QAVaJLdcUh7t1YF5AhPzMSIlK7ul799Xlnbl9VMNXcMMJveB0oaz8YZrbs+cP2IB8xmLJQED2LaCffocyK64GBUVu8HP6bAaiYtYh9WTOUJccOlpUm0K85xq3
RVYHNSdQRLxCuxTMJHS5hfjIJ14SwTfouiBi4iq7IFqf0qfuLLNqFEyxP3Y/UgAxo77RKTf5+2YPc5bh1T5h+GlBy9R0hBGDXT79k2xLJFMzcS3b+1qlCpdOddcELXBA
aZ5jGArPsa+QKivneR/GmefIotnA5nhLmbzVVxvPhGR5kuGBPqMBzvcw2WJkFXOAd9CYwJ1NhYQ43tbz6W0S8womJX6xEpLT3aPHtWJvqEOucEqb0XhIZYX9dymUbmJI
XkrFFBqYiXSfcOmdzynSM7FzGelvp83DNEdOnm3vLwqtXw0/pdqReO/E9gKM60dv/Qo4JFfsW0paTTsyCifkt9zLJnwntEUAmXRT0Z7aXwzmtOhj2SY+AuaW/2ljEsp7
6y1TfGLqFxSO9P4bJZmHMLDqea2v6xUPVma8Fzt9zjnKxbM4orY1If6SeB2C9wjQLd50cE3gDCD9DMmHwcIt0VSbcJUZJeqv6LPJki2nTpAKwTGiebaDPVFDUYlIm2Op
j+LQggWtKyNzhsFCiX2vz3KjnILQmBlSqH7pEmJLQcWcuyn5ttTUsJBJYkPxvCFdKiz5LtIj4P5oR/0Hze5G9Eg3ZTPo/GDb6GC2Tm7XjWxuRz60N7+j7DAvMhBkVFM0
4zIHUle7YiAprA4DepRHPPq6PJ+2heiRwwYSKEbyX66i8lyQVNrVHMJsm9b6/CIzFMezfVirXzAwQQVSbrZjG2spNCCxPRlUHP98UgjM+2HHe46T0HczknoURjzq+N77
2lY0BG0SR4CKf1brIRxK/nEU//VCQRY6DhwKALayqVhgc/hG5dYSOa7Ef3UQZXMGAE4eV8cxnjT3IFpYxkf0tMlpvpxwtgNUF+0GTdFmQWrETliD6qiup51y+Jq7AwiT
g5KAVWnnaCt3xvxhC/Ws4Z/QdwY8LBOFW/GZh5ebzT3gwgxjUcsPFFAGSEFOOJCP961Kjjok0iHYUyDIOR1YrjDDqAmfjK1k2sDcBT9bnQf0QzdR99rmbFuo0t75RSmu
GLkkhJZHtnu+HJ0gRKdI3Fnim7mYhv6pACFaLt19GMDnU89p5fdElSwOIMtKycy3kipe2d6Z8C34mMnQcX9LIoO0UcUYUvfxfoLkWzeI/ABmLKOi0GblAI7UkY1wR2DB
AcTvF8gwooMKmKArv5m08HfXQRzKr5h4dvxJlrcUtzSP0aSJnI2ZnA3eJuPZ1zVRh1E5cTduSpJJBzAccWkBXdhB+dO2xQyVXIq1rOmm5czjBEAvG0Kd4qdHpoAg04HS
4RV5gG0ei3t5gVs7eUGIAXT1zAe574Ks1MJLHI2Haa0O4LnoqsYNqO/z/bXznuusMtJdj1mWFoEmpt0uFRtinH3aU2zVoi6NeEvaFm9aHoN8BzERgy2GofUMEoCzpWjG
G8zznVVaVUSaD/8mwvDgdRmMRaXLy0CQoZzD/jC99h7H1LMXSwCg2/OOxLLAfpnaSDdlM+j8YNvoYLZObteNbLxK57Hc0TjtZayyYk9GKHBOG1yL8mmDS4+xF8ZftoiR
k5nZ5fvexXRFfW+2O/Ra6QHpy/xIFgTodQN86LYc3tb8CvFL9nXrqXZvAioIb0/7Bo6Zhtiml0GC8vXCgccOaY4wUO+TxBggGcuMQEDz7mcyWxNfeHEOxfu1/2FaNJjr
f1XmWeKMuMWfg7yuQhFDZKQtlgvq5Hp/YwOX8NE5+nmmh4aATdNZKofNFJpSQZKRWkhawBopCsyS7G2GQPhHT7tMXcfpQGr2yseNO0ctaLlfG+XUsfkNjIg3lxk/YtGH
RguWJQgUjKP2eLt2XTmJn8qIJtEmvYeBjKtfeWMCbYgsk+gordpNwWyyyukrU3j68b0qqSjGDgcV77iDxmUsdJ0bvupPSkv/bkE9dD0OoHK+mM0b4r0Yxl8ghQ/ZfT9n
chMU8Mp8a/uUUGzAEf1Y+m3yeqr5EH4nLNvHqEHlF/nReobea4V5WWwi8rl/JxixhRpLd2kw+GQIuunn0vHioswH71xp2I6eRNDSVOhy8XogyFNZXO+dhMXr/O3HKCyH
/wCw8Z9KwwNpYlpQeXe/v+Y9wofYoU0er6HUrtwhnRoov3ppLTye9Iv4Vtv/Butmqy4pCDUDcpdPtEZ0lvKMFtynGNtO0SyBEE/lnZbnnwLyrvAb+4wWQHaF+dFO0fjx
yFsTygNU349lzX4Hm0k1Mi85HFWKTEL7+vyb8LuxxrcKkLtdCqlqRjFKsu3HBWP7++pQZWVCU0nEpIMgbRTSn6Net6bSULUZOAw4W9t8hzwL5VryB8pxTn7Fd6CFWpoM
Z1JX8ELk9wDzAHi0BB6ilJWh67ZHT8koe91cMn49Mn3LGtq9ovuKJx1vijJ5gc2eveKmvGfJ3tTGzSi8n2tEzL1Si4IfL77MBYEtwnA8CMscGl++Apc7LV/DvqxAf5bs
7oZar2TcczsftNO2k6tHaX+Sv1M/UJlnyLvRrGKq8Wkdap5WXBOwrzw48X66QAKWcxALD8e73oO9k+fvVp2uPYIeQNgh8mpUkRoqiVFWL0Ut7iy+SKpkpSTvWdC+BjUj
cHPp01BUsLTPRayjhN4cVdlUeoAXpOKRTmIG+zZCtVF9wDEUQu2VfznMy2scSELtXIJcLm1lSxT3cP/gTJIEcoQfdEagFKNR5sYgVz5rreSUDSXaa7JQdBiFeRLpglWM
J1jjWepsd7xC6mUWI+nrwRT+1TjTui98aEHKBNIdUiEXCY0KtcSBtq2tALw5omA2AhRF9BFInuGYnDImb0+QAC4sIFovItFZuV/UjqgYVqPrK63Cu6isTPIDjccXUp+c
hB8/T0FlP/gm1KUNBLWexkVSM4IeRY91j2vionTwoAaQh9zOQnHKfFCybvkFyjtcsUdQnS2NaP2sJWpX/no0fv0bGr+3Vx0Rvts2vtp9za6MpQkqhXzR3m6z5QO5HMlB
eUS65PDnFuugIkAARwxu2BNNwpu5In1wNPj1bx8tzVQY3NFjY4VxxkltajDNOhpvPduiAujzgeyRjwj8gj3DM3gzsgjR+uAt/VwXWVAkDF4YCet/Up8wCKNUIfuvmxNW
gB1pRi2Y2eGdPeS4k4N1IZFy9EJsXfhoGehuK13C8pMIBZsPijDxLcSMOFX6/G8WOyeu7JN8lsK0H5GdduMr9dx9ocVz+K6ZQ0JcP/YPgj8FovkNHWgCsSGCMOfnFHMG
7wOyRKukP/89tAN0xm6TXwz8InDPCgHgk3K12GRO97mn2Q+pGyOSaqRkbBRWnOlkx8im485+tmWiy8ctb14yOJRlPm8K4Fx/RcQj8V77HPoMWacmhheSe+R4gykAUMcx
Nm800/jxXMweIIZMWcOMZ9IVrolBWmxKb5b7G+3uF4WlT2Mbaz5BAbqTS0z4aLSnGWqVf+/+Fiv1W6RRP+0eG+MY3iwQDp8Lqr2t5cfdw3POaEdiNitYss7kQelk9ERe
pDgzMi/17t80XMRXrkwSjH0MFlno0iSfkp0uze9bUBAfWEY0ZQA2wHDUjKbTaZke9aVwqvfAnc5Bl3h7i1k2tc3bNu0gJLss+nJjcYhLwlemkFykSinXKRPG9GW6/UP0
Uu7B73QIikzIEvN1L9W/qKFmcVhNEHBcrmL+qvRiiRXbRbGqZgBIZmRzIfIGY/Ll4MIMY1HLDxRQBkhBTjiQj8KceLc/lUm8SDMDYD4RJYeJjACH9vBU/l5L033Et+YM
ItWxMHGXS6d4ZmHeyKYpesvMNit27U+QOs+hhAwrqT/8JPg/9fVH0FcIplyJBK87UZvK+VYsgFAJUup7xeOT4yLVsTBxl0uneGZh3simKXqbBKKQwWJwHz8mOdF3RUY8
YgSKxTItS3FnWW19ZJdu3I9SJEUwD6mPKI3g4DdWS+1gqcaGWATF8OqGxohLG3pajHgZSTvNKAmLy41G5rDlU4tlG5Ew0kEi1HUSNFn6amSbGdFS1EE6wCQY9zv6+ZcG
8ckrJD1fsePFDMdxBG6sIyeoXiRoMeRXuaIzTADEN4IK+9Az9FTTq9tyq0wu+7Wu9xL4yw4Fnwvb7Z8n2tCZCFdvCynfbRwgbvqdNR+ACvLy7chiyKTFrGBqZTvJ2TQC
kBHYubzzrcSO1O11GmPNlS93zE45n6kKUV0frtnVhv0dq8mpfABxDKm7zfTl9RHhbuaWGVYEvBtpeBUv3akNhgtDP2YDexJbofrIGOgqiLzyds9TQhryHA0lp59Z8vHA
fax7nH6nftQkevEzKJ6QuYmgyXG40Ofsia/OO6Y7i3jXTHMLzNiFb5Y51Z6IZsTMJgEn28BD/gtKU8qdGKySviEHN53mfRGwMsVLyIRFfReusbcIwP+Dg3Eyr+I9oKjf
HavJqXwAcQypu8305fUR4SFezK64zQQHiDaQRlynWUouDpFXuAp//waewqHLejtvJ6heJGgx5Fe5ojNMAMQ3ghiImNR3p0quPT3ndUPJnyivVkwmg/osVBBhNEie+l5l
ulfVOwQghnrZBOFIqdXwaZOjnZNb0nEEgN2pCilQzz0DMQRxChpuYtJH9GY7NkkS+CUhZh7jMPhYUzQatmF1dCYBJ9vAQ/4LSlPKnRiskr7tQKevc8fpYjvKD9rjnUoe
2fY2VSUkfpTZjSgdDaAwHt+VtWEEmx9l2CqDSRWZ2NYmw0u+CoL0kFWpu9gNaMllnCJQ/XRcLSsuBqiIRH8yo0PsNNTiSXyodTeS0AeuvNgR9xrPrkD0XVyJAWYxsAbE
ZyOf+F2Ojrxj+H1oaVo4fFYBu5q6SDJs5mjfte2eCod9Ps/N1O80EYkNMATaMSIbhfiSyEJVMk/nqfVOA9HTySb44RazEyaZFkxhWuxCZDx7D3so3pYqivzrjZI2lTer
9M1/YPaxHUyFmifkeJOET5hb1XYGpH/W90fsNYSVm+2Nv5Ee3NDXtxi4NElH705kNleuka9udbk9pZPyQ97Zx8fLUYQlZ9svahLaGW+8W4OE13CJI4f+NXp3CCfb/z3D
awbE0ZQ5A5lQrc5BT8VOE2cjn/hdjo68Y/h9aGlaOHyQ+JY4SbAmfRzS9zR75NwCfqXpAg7kFALpeRk1yhJ1i36YivpufBI5UwZOPm+AeRaaoqBs8Gu/KcHj7QW3+2Go
O3GsTLlJVbJtE6RXdxgCfEg3ZTPo/GDb6GC2Tm7XjWwIpDSx6b0SYweqhQNBPuIW/Fp9zhBqVYGhekmXj4s4WuRKmve6sjJfW2RjjCQWnakTpriKnsS4lKig5PJ6SwCG
tydAnOQ8tCFUq7qC+E0t07k60SibFvgPjefwCV6cc9ArfLIFkfuf4uDxgnOae69cz1X+pb4x9iKokSGP40aE2NjS9lAHXWCNZ618bOMvghofrG3IbyRt5/eRtdJRzNf4
ejobVQ/GGJiJEhovtDILFmU21gIp7b4nZrsRpkyfIYL/qpyNnTv6rt/mYyfMTYoP42c3A1jQJsFWgTkIFns2tJskV2lMD4/bT+rqVAd74gdIim4a+q1AD5KHUn90lqSu
QajWoqraTlYyh1Oh22I1Atx6tydsF372/idpOww1B5nY0vZQB11gjWetfGzjL4IatrA4g+RJUl3qkYLWdaEYcXSErWzJ44Mt3+aL9xFbbwz8Wn3OEGpVgaF6SZePizha
Ny1CdLpQ9iprrMptZywASHxxsywiyB89E4j9Ac4w22RLXvJaLjMr22ADXB8Uk3mHcqQFhJFGmcLmP5mxobupNTMNFT0ULwZF5/gImAqRIF1/sioFgDHmp6jz8bfui46v
SIpuGvqtQA+Sh1J/dJakrgNlJBGnj6sjYg4h57MHymc279faPrMA24ehCwqcIgsClYx6sSB2RmpBE8PKadgsvTbPlWEY9LyY5vK3BOKIBQcTnXKY4myFzdJ5zJYFjsy4
cVOJe9S5JfRH1w9Ao9dSz+LD0J/OcUJ6Y8I0Y2FQ+//8CvFL9nXrqXZvAioIb0/7ub9ln8Ysl2W8jel8lmYAEARogtVO4yTrm2hzurVhJzozm+ZkUNdQWxYUBo5J3IJg
wpx4tz+VSbxIMwNgPhElh/o0YZ9cTYOG2N2GkI/drRRGLQh9hqCEjlUrk9eTS+NF7JPR9+hzQ1ticbKVG+Y9svetSo46JNIh2FMgyDkdWK7Vi9Hf4HRg8WL15JsjSGW5
bEtsvZDRkUpbQWkWDv/V1CV8TehI2ZCZuvIL1/pA2mV65izJGiMSr/wMXYLJH/5JNYC6l/FgUt8Zc0TKd8BA9pwaKhz+qzHMlDLbrZ2M4DQYQPTAI6ugVkb3UlqlOlIc
SGYr4zikbOZfwPeZ0S3J0uwROQBd4izSzJaFpiES1zhDa2o3T19BPi5rJr5UJLHsYsHLt9K7DUim4tRUQqlPgKQ4MzIv9e7fNFzEV65MEox9DBZZ6NIkn5KdLs3vW1AQ
H1hGNGUANsBw1Iym02mZHtwrU+Ndw19dxv9dv8HjP8QpjvxvDjbESAEH12N4m7C2odhHfprCfygemARTrLHNJ7+/6nT05GZRUkKVyyjyI246p6m4Ml53XwwPVttl7Gly
g+7W7ZQM9KMjtF9YZ8aRy/ETuDD8pqq8Bb1PNa1KhhQpjvxvDjbESAEH12N4m7C2odhHfprCfygemARTrLHNJ7+/6nT05GZRUkKVyyjyI27JXW9j4sHiXWl/F7zPC7Tc
YgSKxTItS3FnWW19ZJdu3I9SJEUwD6mPKI3g4DdWS+3eIW6iW1nXAc/op/hFJ23VjHgZSTvNKAmLy41G5rDlU4tlG5Ew0kEi1HUSNFn6amSK82GKLVtZRcHFDgxoVK8+
uD8cwAiyPTaD+4ObMHiFsouGXeyVOVpM2MaOxhYJ3VqWWi3m3Ltzi2X7Wg6ycd6FIS8KoO6re6/F6dt+Ln6wK4ZrpcZHaGmXmVwwHwomqAkPC6KzbkIromz2J0Ipocmx
gqpNP0dWBizTO3FEK69tsWk50iUimmmW3gVZs0NvUfS0lEmxcyVz4W4tM7allcq/6qujaX7J9Iqi5auzfNLa5DLkXLMl+BDGrwcAhElGG0JwulLGbxYXtdszLqVcV1kg
brH8xQLaoKG9COvwikTRnGhhL78a2VICVwR8OjiVaF3WriYfBXbOQIqjZD7sI0S3U8wo4ltu/ZJLah1J96j+ZuApWpetS8lSFC7aqdfbFpj1SYctbY/1kT0CnyGgfQUU
tJRJsXMlc+FuLTO2pZXKv6XAOgDekCZqtPUQQfjBQJ+wDIQhp1zNmrCpMPmlx0uNi4Zd7JU5WkzYxo7GFgndWkqF1cLPXmtXntK7wyBUfAAA4Xb9V1rceUXS+hj4UqNx
NEgb2SBD1cFPLYSq+QnihX+xBmhVngfTW0gJAIAYifC9vfkmLoJqQZ2AZ2Ft8YwbNUbeixYYzOH4ORv7qgUwOlPMKOJbbv2SS2odSfeo/mZQgBx3u8PChkMbCB0Y4aNU
CsNVoCISRRIgzeKIesfCUwvyKrcBoeh98CI2Qg3cggI2z5VhGPS8mObytwTiiAUHE51ymOJshc3SecyWBY7MuHFTiXvUuSX0R9cPQKPXUs/iw9CfznFCemPCNGNhUPv/
/ArxS/Z166l2bwIqCG9P+xnVDtIvGyxv6wwXrcORscoRhq3edEcxkW1mmKZBYrxA6n/ftlsA850SRmz+cQSLoNVVgdoFWgx/fZR/C3LQHMLtdMiPzawb8vy7rjv6BZhp
g+7W7ZQM9KMjtF9YZ8aRy/ETuDD8pqq8Bb1PNa1KhhQpjvxvDjbESAEH12N4m7C2odhHfprCfygemARTrLHNJ1nnLnk0YI0G8DwUQrZUmf7sETkAXeIs0syWhaYhEtc4
V6gkWfjOoEpiQyhLi3XG0cVoDcOftmJSkNBRohfQY2n581x/Hs+drj3702OOnUMXGr6rM/CxwuXoNMGTf6nbbKxVhYyhrteTNFcvZ51iXwJX3jzdKhYMF4s1ODZ5c4Oo
1VWB2gVaDH99lH8LctAcwmwgcuKpVOD2wRb+9zmQbxkLQnSNCohHvPZezIAyyoFe0d3ic4Qavzqocec4a1eSvwuDp1sUAbaM5TpIZhp0vzoWS5vIP0RT2SQXsmc2eu5S
PAB2/kNlWR12cUMBTmPU1mR3yZ1AJ+aGbrAc11Jgy1f7ZeSm9g9X5vWkKvDJStDI0PiMkdfnJo+WIpaEIr0goHv++pkOUs+k1XcAtFLMXsOg1v1jRvfXgbT5zLj1vfkB
KY78bw42xEgBB9djeJuwtqHYR36awn8oHpgEU6yxzSejrblSOvyLQWAn28PzXVDis/lb+RisBtnq1hzpEKVmtvG9Kqkoxg4HFe+4g8ZlLHSdG77qT0pL/25BPXQ9DqBy
fLHa1OcVXuzZbfZTj6Uvs6B0qUHF4Mv326X3Gx7iDxHPHyE8HNbEyjrcR3P86La28yybqd8f9mfsY3cspq1xBOiy7g009t8vWqvxsEdxibNogzuuARDz+fqqmKp6K1L0
5rSY+jBTGZ35Dgw0GxpEBpJpR1uPFSeHDIA/PXhQgzsQVYpg8jfFkpQZMAWK4dPRrhskJafPL4mIFo+zKedCkVIp4JzFNe8fm8nYdIUNOaeYWeOX/X7NNSs1wGg7jRhg
0s5E8+YOAU/H61w1ewBE86fHHHd1kaH+2ssrzP6NwslLdC9q6Z0ysbqhU/LB57ag554MO5kscjzWvYIN6aKcKWqiZ9t1tuuv9up4gRaiPtUPEWaBMozMC7en1Eu1dn0N
aIM7rgEQ8/n6qpiqeitS9D/I1LWMLvHhKHnmzIPpdQev6gdz94CKgxE4GzEiIf3c5XUO20fHpn/ZZM+rJtx/EzRrT4YXOmV8RnzSM8KOQe/6vPsBaDXQvgn1uIsV5QjY
cnDxWPaILTh8fM/7FSib6cv4KUpRfP/E0GRMNmnnbHJpsFlAVk46VVAlMgI2vSXlo9H+1bdD24mRK3hCloZI1Hk7Z7ZXtVdOZljwlBKFqhaE9xYBsaHENJpoqHo5f8G4
4xtqAF+++AefGnMPpjS2Q3hcGl8ImSJP8qDDE0sfOq2sZeArS+pMcDaFB9saMHJUiY9DbwBJ1/5LaSlwUDuu50HZMg9NXGoKyOp8NrXMJPLlm7kc+eIxjHB2DPsT2Ed7
79aQ5j/Bnl8ltfsJgIaX2O3RfO0gooYq2UZ+fmTlALkv0mKUlp8Pp24m1H6i4ZV5yT8HCTawmc3euzXYSuSUi3zY5C87A5cp3khR5gjfKKzqM3XxhTmznePOpU4FSDCQ
/DmAbsSiKI+XMPCyJp7/m4mPQ28ASdf+S2kpcFA7rucsG/CIj+/mMW5KWTrBSpe7azMSuIUrMZRtx9uBaJ6zE2mwWUBWTjpVUCUyAja9JeXU2ytvg+3h6VyfsFUOr7c4
oSWZRl3aEO3jcW+AhBeb5edGUx5xYVJ+inB3VFhdAM7Cdb9yN/RASEx4ScG4oThxOm8JSebrCjHzcnlyEWAWwSPCtAkzJTCvLOiN23hHLql82OQvOwOXKd5IUeYI3yis
+YgM2K+Q1n1ajNHh4b2wFaLQEhoMHrdKFWdJNfo9MUt6fJNSxmPeVwggWCxcKweBj0lCmsAMAt8wG6lzQSRBbY4SkDINbxogquKyngu7z7Ii1ZoQSBS4/WIB40qR1cho
G585PVlNi2E9TosT0fmx3DMiK/wnSe6YPmXp+I1w+Xcd55SvAgULfVQKteITpIJr0pFiezxtXin6+Fyc6DDJvkwQDevbANLdFM8Towjo1c2+mwbtA0ObMWpWXPBwFgUE
xKCLppop1BYYZIF+DUrXMa7ul+9fHIGPQo8uY3s/YosvgQKLU4h8B/oWbt+TvKx4X/hKANoXUAPFrssFdhN8vMpT36fgUaNoO3gq31lVX1JXLBIB2dBFAKgiGpD1PN5s
KAUddGqzNZrX/WtQxR6MxOBwNr9RgJYv9cj6mzml9ZqF7llfJ22JqbVxGPa+FM/ff+0fNYrdN8uyGAPqpumO551kCtoMlCsbC9nc64s907gi7s94rTCq5MV61yBm/8ov
pBlvJJlSVH5o09J6cNfkHxc2DodID6h2ZrIPh6l7ujUJU7ZyYgp2tRuZXmKIj5sVysqOJzg0onpBmyJn4V8xOyMSsR+J4NMinIU4uRD0LHRjwztQKyz+8mgShtQBNnMM
vsW5kfrNCNenQLpYAwyePKWPH1CHRG6N7z8yeTVAqx59w1p99zxCEL6rCuX7rXTLZhq3zJn3psAxOKuUBwsUqlCLnLTYHoK8nhL5/rXxQuJxBc5+r3DodYVSNz2+6kSc
rDR7eaqRQUV6OKO/1VvfxsljKFAR2Jc5ZrMHkt2yePQzRSXWzyQMNgT51L5F7CnUMI0OzfRHFPHp5Z2w2PWCtSGlOMLqTsvj3bP3p1Qt0jTWJ/suScrSNGaFyyl+lyoJ
/xw7rBuetkAN/J7cNiDOCnJw8Vj2iC04fHzP+xUom+lbkp+9KQbHQm69Ax4S7fZi+EpcNXMxRmp01rkIzFw2FoOqNeTpIGRqjOycBTuIqnOshU2ty8dqNk30SbiOqwv5
+2ZZkgJ6RGIwbM/quyqy6xmOO8mY9Vt21GWF+tBZ4jev4d1g0OlMLEK4W7lWHCb2zk61/796DMQSnhkr6GunuegKcnRunRDW5I02sjBp9KiObaNFT2vmMvMjGJ1D/8BV
Od6LMeGFSNlt8kFC4PlKNhj+uJL+zKrchZaef9gcOT7tVv7XmNW3zwnf4CrlS8MQqrfxEGqeTW/F2N/HZq0I33HpPUW36qcxgw7CrT0NvewwzUV/mn9+QWeqbyNtKaMO
xCtLTaJb572inH8IfjBU/rTLpAp8V1UHiK0MZTKvhX5+rGfK/+Fiw5v2vOSJGowDAtyej/YrPa1np57jlMPHVZXDCJozNsicZI1nAcV10tU1KMVWZBBqU0epGKJ9CNI8
Sm4kKsGKLJEwuMcKy2D5pryZyKIBNqJXaXFH3Yx/cGuL50Mxmt824ehhqeBUcZRzZvehPPzjvxAmn04UJ1Vf/M/Sudo8q/T2PTGPmcS/go6QCpqqNEtuxXq8rpFTfSQC
O+HrfeDfY1OnXZQnawneGJ+uIR/boAlg2tRSee2i1amLVmyZ3vtpWhaq8rkTIF+54FYJm/PqkaapdPuFv4moVSjwAfDj6tU9Zmm6YHy3AU9rzeSnXLGvOiQkEp6unbJ8
4KujpQREnF1GKF6LuVm9m7h9K/7Jr32gvRw181tMtBZhumcrz2wS5AexXaUo9PL68GFb6UC+yi+y/lVda85aKdKrrFvCiVDqopqOPfb8D2C4fSv+ya99oL0cNfNbTLQW
YbpnK89sEuQHsV2lKPTy+vBhW+lAvsovsv5VXWvOWimQH2s3smFP7KMOUBT17QZdndNsfA/1tbJgPDBRsXFG60f+tutYa0YFRilMUCa2GwhM5Nfh8dxy4UJp9w0x/WoG
uJSllM3z/+zPswBNHII8r2tJET244Crm50XAm2AUh6HQqOTCpW6FZUSFjwrGoMwAaI440oaWe8aRMsDM/iRYCeQ+qPJTlQio3Crpg/ZHrrd14VS5C/zR9/F5zTQmZxbP
BCcTzdXqNApimHS8tKeoYmb3oTz8478QJp9OFCdVX/zP0rnaPKv09j0xj5nEv4KOvn2ASIi8EI66gDyA2XAxEx057H7XiWh7K9xKdwV86YfxYalwBnUdqaYzUwH1541z
+wSGJP4JCzIu3pUAEL3wjhnIdLjxc0AckyP3Z4CNe7MwElZwAgjBan9CuDdpho34fw7L3OlJXtAeZBNwTotiUmFUIgay7Wrn/kYlVNX4qZ6ORwen15l47gBfpxVN0LuI
15fJcjW7KTY3yDaZf2e45Gm2J6Kqosni0JgodfpGejS1weazumorvwETrWLgsljlZguNhRQXSvjqkJzzEzkT4svsFOUFzdHAiL/jFjmHJNGLVmyZ3vtpWhaq8rkTIF+5
4FYJm/PqkaapdPuFv4moVS3AnE2CnxsLoY3prfc0ITfxS+KgOlPONpuN/a0vAp6U8N1aPxmevwymdDSlfwHvUP+8Xo30h+J03kpgzFz58YCuhYu61msoBRfZlualkmyk
TLRCclDQll95i3p5mTlhNnGRw/wt0MGLicNTyaXRtyvCNMu+qm1toc4FMKNGthR8g0hb0XqzREKVqWSo6DgCqnyRRsf5IgXQbZMvXiuaNJGl1C/Af8aKGahJeK9y2KTX
CYz5N0mcSa1CzgmYXzPKsrV043iO25eP5tzmMEcnapbL7BTlBc3RwIi/4xY5hyTRi1Zsmd77aVoWqvK5EyBfueBWCZvz6pGmqXT7hb+JqFXzzEHOuG6r7yuw745fJ5TY
Gf/DFYSUkceNiruL1dNbx8NDKsvzx6+MmT1Qcl/4dXeQ7UC2qD3lKTe6uOu0/TfTRhwiYFxo7k/2bEgcTYAVNmDkrGm6bEGlNlVflRgXHznVKZdbnbHSvEBrq7qIh5i7
oOnLowbvOBJ3ADyoqd/KtQhfpMEPMK02oWq55fP+pFeWnTJr/9PfS2jsaIIAZ93VQ+w01OJJfKh1N5LQB6682HFachhE8w26Wr568IjO6jvxYalwBnUdqaYzUwH1541z
2GsTZa0bvSd0dYgnaF6MgIBsxzqzhALRgye8u3ucAnlhVCIGsu1q5/5GJVTV+KmejkcHp9eZeO4AX6cVTdC7iPqpD64ZeYkulSXO7bA/4Sha1fV5Kdl7gZHTafmAjO1B
v2yog+W/vKV4tpANrZwVtSA3XWSiOEwWr3SeLxo582+NajTDQFtyaE/9+CRPp/4huH0r/smvfaC9HDXzW0y0FmG6ZyvPbBLkB7FdpSj08voXwuWhpJhIDBDsFyYcCsb8
wqgKhKx1HIcULS4g3iB36jqjknTRWQdquVBNQkW9bs0tLDoSO3SwfaJU0ma7tbMbyDbQhlVsr4GWGYK+bY/Zi8I0y76qbW2hzgUwo0a2FHyDSFvRerNEQpWpZKjoOAKq
r2qC8Gkq9aEpiM+QZG+M9hOAwQNBTwe3u8Dum38iMuKqZgf1Sru0vgMtJIeqEpMb0uwar8UbzPPHVEUG8CvD6dYJ5UPb5CrDQRbD+Vt6RTxrJDURTMeQFoXZ/TeccdxM
eWiWqwzkUedzd2a6+vgBUhiKhxrb5Voy9fSfi+Fl3NJUu04FIU9O5JVK5YTndFXi9EQYRGy4L7Rv5MRtbsmV/e6BjvaHy3qbc/nHl9+x785yE9AMdO02tnF4mE/RaXkC
kj4FKZNXJ7AY6jwNJB07PKBA8/Ho5IJHGXIlSW1V57tCxjAm9qycQ0B3PxhFh1peroWLutZrKAUX2ZbmpZJspEy0QnJQ0JZfeYt6eZk5YTZxtOWWwk75g5g/bTAshdBS
Gf/DFYSUkceNiruL1dNbx6fXRzEhzrnpwvYZUH0sgt5vYVuIFB4m8EYD/fWvI4o+L8IqiTNs7v7I7gUquAXd00uzp2VkwGZ3/HVjUp6SuAKEdJGz3kB1U4BPH3qpS3S6
vJ94oFL04Cava73EnEdNDmd1SSl3itQ5p+c7xfNf+HzH1LMXSwCg2/OOxLLAfpna6ApydG6dENbkjTayMGn0qCTJxpuh9tdKyE7+gvcNUXNc/G+8T9WYw6mynBo4Ye/6
VLtOBSFPTuSVSuWE53RV4vREGERsuC+0b+TEbW7Jlf1p+FUDEXyZSiBN3wiGnggfOuFwFbxVcgr7gQQ7mFvRzsjhYp+LITNIrLVY/j1Da8QdX8xHSb/qAKwUtZR11BYf
hHSRs95AdVOATx96qUt0uryfeKBS9OAmr2u9xJxHTQ5e9RmaaNhxaguVJGCiNMefOuFwFbxVcgr7gQQ7mFvRzsjhYp+LITNIrLVY/j1Da8TgfwyVI3l1ZksAwqd9v7CU
hHSRs95AdVOATx96qUt0uryfeKBS9OAmr2u9xJxHTQ7a06MH0O0Kw1DI/BieNVzcB1Rsg9Wea15vJHZCu9K4tWBEHbJ+aytYHbOH4zLkQv9n2sQ1IlW6xYChbzEqtyoi
S4f7+/7ddbd5KEX/ozG2zMsKGI+e2g2S+8TaQyydBZvJ525uvIPFFBIHEk+pgKNv6ApydG6dENbkjTayMGn0qAYwc546PUCbMF80PxTE20pm96E8/OO/ECafThQnVV/8
z9K52jyr9PY9MY+ZxL+CjuT/Qn/CBO2Pn9KEVEh7Q8VK9nQLAZ96bZXY1nRubCwTKMaQIL9FAyh2ocUc6vGSEyvVKylVQpOTEtTmJc+1s9JETdCG6JyI2aMa34YugmMp
HWeIPNSJPn37ryisqxOA8B5r1r3g7//0f6/MbWe5YDhOuERHHuZyER00TKlOjUxWZ/lyYc5uX9FLwA2b2waAI0JMz3jW2JY+iF+BVT2k6JAjqOVw/CfWoMONZe3mmVZ6
5dqij41m5+rsOTQ1uparYa7ul+9fHIGPQo8uY3s/Yov0YRimBllRFRBHq57Hj+qnBCcTzdXqNApimHS8tKeoYsf5/wSkKLdcmpMLEUoqYJ8SoqhpFTy9bB9JYLdaphCw
8taqJXue+34RL80Lj5h+OqHQ8Lb/521rhjLoVMECBxlkHHxCajLMldRi9HBYKq5OwtUfmSULuE9If2FSGZwqrZ+AUxHdCb71wlx73LaEYCi8k8pKiPwz9dHP40evHscT
/c7WUfu4ioEZ3Gxg+HkKR4tWbJne+2laFqryuRMgX7ngVgmb8+qRpql0+4W/iahVwP1mYsURq2Nv0FXeigvC0QGiNtbIpIbBeGbfbid/kxrVKZdbnbHSvEBrq7qIh5i7
nkEeJWbhXsFT7wK+c31lm6UVBhV9ewOed/Mvc5OHtdM4zDN605iltU4yycKNT/nQO9dlglVwxFM3K97yTfzN6/29CWnvQJjzmBf7ELLbRd5odJxjcGOK7QHrCpXhRWQt
RUVp4dcA/Y0fdoDZ5Dp69tmq7IBBBThbX48YIRRHVXSzPNrcS6g3UliuSsyeYVAkp4dLWCW+eScEndM7iVU+sQ2D6Q01zl0CHT4qZznO2qJs/5qntXMOjKvHDry9weVM
zKw91Zchd9ucxO5mTFxHHfX4UdfIlIQEKjGxeSnCI/B0lPlVbrADNbJ7iNb/q6laQkzPeNbYlj6IX4FVPaTokPLWqiV7nvt+ES/NC4+Yfjr6qTwD6uITDIy4mE3GdIwa
nvUm4OWaNpBPRoZ8dPRlp7RNPZSY2tVbJl9SrmWnqpfXfwmavFUpEoZQfYCyzAS6XsBRfcABy9qow49SBO2iCGuJ80SZzkey0yqvkXHmKQ8WE7yJVU3Fura1OJm+mj27
cTcCaT036ITe1kKmIMq6TUN2+mdVY43DgeGvHCviGAHvxYb6v85XaNRq1clLeo33jWo0w0BbcmhP/fgkT6f+IfBmIxMdnNWtkyXd/rsLrCr0lc7StiSpvdCaYDadBrpa
YVQiBrLtauf+RiVU1fipnjRk3rS3dX32gk04Q8NVTSWHClFfJUQ0Yln9V55VJydDAHJgYnetRbFIpFaSqRNcGjDNOswLA9rSdRp+HZAEsDbmiTFU8RDyPNzZCB+J3gvH
e5et+oAKNUPhIHGTmLyMFK3+yn+d7JU5sOOfFtfFu73SaolOoZnRN4CmSQPsQ8QdiD1oCYGkyatCb1d3g0apf38Oy9zpSV7QHmQTcE6LYlLjs95pBtU2cBp5E04dZQW3
ZvehPPzjvxAmn04UJ1Vf/M/Sudo8q/T2PTGPmcS/go7YD8g6QD+m0pcGkjN99qN8uUmf74jaevfgJQPE3/ftu9d/CZq8VSkShlB9gLLMBLoEsv5GjSuya9cW/dUKeBNK
C3p6NymCjzkZQRHJtPgSfDjgGQAfwUgL14MLQ5eind6Zh66GAUlIjTo3EFod6u96JsB/US1aiA2AuwYP+beG6Qmn+N1vNrAix3SEsiV9pz6BxP+BwMsHPKxhxLbF1Wg1
dtSwmRK7t5DXx9ksH/imYYtMIj1E7Duf3ctXt6qtHOVi9CGUKwBAvXRpuPn6UblAvOWA9vPYxdak/wp61srTU/4ZJkVkpRTcCUVMvzLdGIdiBIrFMi1LcWdZbX1kl27c
BbZO5bvudqwxgk3+WcrTxQQnE83V6jQKYph0vLSnqGL3dpwKNCmryKWeQR5dyA4YEEHbK2RONQ7likaebCYPI5Ljm0kQiZ92+jcEsEco62VqayJC6guQaPFK2TSrDTuz
5dCPxfDzS3HFeh+jjfcYcdv2yrZbIQCHY3y8nboRbUZfYzzkrDM3HkNXFCxOHDPNn/lBtb2T9o1s6WwMFfBZCQa82JN5LIIJO19G7FJms3FibuDieN6/6YLGJ2h3d8yS
Z2aANdrCFXBQQSauB2fHfUsiLt+a8sSjtJu43cym9C715eltlPUWMD/JFxAsynZZqW9esK5c4Fwb3KQBdOCeX6BoVCOp2OHpwdg4S88+7JUZOr0GpwSqtIKrB4QwcYzt
9UwHSRA00kIh99vyFVHaG2nXlaxhD5JENJuvvbD3yNlgE3kN1WwN+rbWRNSijf3dQMR4TZouJJF7lo9DVsXTvykZpRaEo2S3NbNhztSaGwZoDSEsqJt5ACML0A3vQh2N
eYNV6wWtjRZ5kZqIsRQyKVSmeGdS0oeeXEwg+vV1MRQJm8zxMW4UKQIE0Yv0qo8gu+3hM8vxRYeAmzB+Hc4V84v+jPE3k/zFOUHQtP4lUJ2HOEJ06e1uin+wz7MWFs8y
UMcFEoZuyy5fEXG4Dwhz5ul1mLujyiVMIEl68WjLcq6AOj5ZRu6QuviqVqVhSVks8pFckG9akA/ybls/ec9WbJ/fI6iWeEK1bmupzpjd38ItzYmOMBL8Dy+Rf8imCddO
hcozMiTpcZ3lqpKIeWYw0wk6sFIbiJcPGhvKBy0oj+rsRc4a7+Py8x6d94jcATROQ2unxBk1az1QSLmPoy2DNDbTeAcYoPfYlcbirQK8/fBXOaHgb2d+wt8/VHRGjHIH
Hj7zMFWYg9ti4FOTSZiZpov+jPE3k/zFOUHQtP4lUJ1y6l2A1of+FKi3ezVvA0YCHVIdT389dhpEgFo96O2xj2nXlaxhD5JENJuvvbD3yNnBzrMKkPfdOAZmIQmAqb0l
36Eg6yyvMgz55vwasoxtLKS0PE42MVmBKCD2jOUzPSsHWjL51fFykTM9QDiQ2QMZSkOrELeN3gPYG4U1CyOK5MN95tSwEWhCRpX/szdVw4yVkYJpIJ1grmilEogVQ1Pe
7UBMsqVRg1xEIh4albaQKUhoqADwFXxAj8BqwEg/kRw/fvkChriLGg+QfiF33Wd9jPkI8+dQkNMub+RoYvhD2gSI9wOvYVUWF4/0SfVT9DLqfPNaMHhV1OpoXVZtchT6
pmwUIpwEyviFRNSSyG6q60PiIDD573fP4YbxqoJgYOywl2OiDNm+qLGP/z1b+pElhaLj7Rl4Q63AaAhIVY1kGKtKHy9XDjN3KIZDJTWW3kau2W7XPMtMOsVPue4apq2v
B0k5ozv3AzciT3JEKSJ2T4nc+cW4JAqVxIct5Zb7IsRkZyJ7pQJFsmxpwi/0djDNWstL0E20RPCDsVYjBWu7uOv8b9ZYgxnekj6MtmCDLffUQDv4w9GTG2i4SgwPoltW
+pQNVTtp1593dl9fZvFlosZO3klobdqbmXXeHcDptSVGdu/Zq20imM2kp3j0QY7pNtN4Bxig99iVxuKtArz98ORNEojY1vofhSonj++haaoZ0LfSgclURtIvtyFwQLu+
fdpTbNWiLo14S9oWb1oeg7rRQfzxktIcVmiSXiwFdfa6DVIjaAxgiHjDfTX1eQYrw6FN/vObyB/SWZeGiR0arMhMmCqSqV4QTQHGmaVt9bgQVDFqWFUGJnlHtT35Zktq
Hj7zMFWYg9ti4FOTSZiZpov+jPE3k/zFOUHQtP4lUJ1y6l2A1of+FKi3ezVvA0YC5j3Ch9ihTR6vodSu3CGdGj5d+MM9gzbljTpkRsG8HqeOz7MC+33zCj+KpP98lWZH
MNgOjhF/zBVFS0oj6q1COpyftzRGPB1tOEqM0UyTtkLPqmjn1lzKgfuh+7aofuKqpmwUIpwEyviFRNSSyG6q60PiIDD573fP4YbxqoJgYOxhs4zVLaWtfsWfCheUBFUJ
tagWzPztlZMWdmiaKMub7ewd4DYsJmDyDNvv8Kzz4wNkZRQmShbqzrD51uvdJALZ/5q2bCoyrND3UFoYso5/dmFLF7UqplXE8p+f2Xu/STMw2A6OEX/MFUVLSiPqrUI6
S1w1mNdvOSG7TEik7Mno0/ieMMy/4XH17Cvs99dKLS6VpVKx3ImLXpZdwpls2CJ3dhw4vpgmV75RZAY7U+XcNoXKMzIk6XGd5aqSiHlmMNOhRJ0meFV+MrD/7rqdd/S4
uKq0GQ3MFrow3LsEfhVKFcPm+BgYdVcMqtepLkN7UuZ39jsAFc5TaXjscGVsJ+7j8gEnhi/MWu8fa5c8Z03NMib6cJ6w/xeyzYwST+kwq9S2STT7fAPOoLBB++3VBSII
fcTRKyN1UTeV+rJB5dkYKQrLx770rcdK7YlPpqOC5HEhc2W/Q6vUkbE2o5oa36EU7TxVqkJWGa+BXCuE35F/x+1ATLKlUYNcRCIeGpW2kCnAsDZC6i6XQevrx+/JGdKH
zsaX973t+w3ybNGI/PqDUXq2jHqek+fokHjWWPSjMrvQxI/OvcxeazATqf2OaqbT8yybqd8f9mfsY3cspq1xBC/3iRpFlj4Z1eu7fngN9sjg2tWkR9CPdT5jTJTcaPi6
Db2NJcbpu1JPHiJ+uGNDYamE3xFRKL5xe5vg8Zj8FhN99dcPt6tsxdtAox8MfVutz7E+dIlB4EGULSPL8Tn/n5b4UQlgx2AN9VvHfs3egNjJAF8x8wdr/E7p72bDZc+/
c+K/Ez3KrtrHtzf1M/QFsbpu/Fmdfidw3Wsbn90D97ll6HlCc9RhDfCCp/ZUNcBVsXgdWmARIacxWQXjUSwxyY4LzwAFl/1TNGWdpRt0dRc842PzWtPDQSIdDlBvPMcY
Cy/L/AzRBqCQr0EBydANvVUjqoUHiwPj73qU/BvL5zOuHankI4ZqbkOwattknzMUhLrKkyKA0FPl+PQC3p9Z0n8Oy9zpSV7QHmQTcE6LYlIJw718ZIChW4TeZKva37tI
bvVRKOCo4fpic66v6ObayJnXxBdvMhJuc65Jmm1uxumMFMFp9m8Fkozjo4hbi5DTiy7s2mbo/n4I76A8VdBP9cYuERN90t+TDEv3a3jwYS+soy9A/pTRFK2jOM+edlLB
Z6jHHAR/fkzlK7ZrIa7ltv8SlWba3mkMf7Qppcwuil0bhS7hAVQstEe4ZhHa1NcAfJdHwq6PgbgQavQXhseQ8Id4O33clQo95Vd4q6/vbJcUwtP2OQbr7jUnCm9oUJkZ
YqtMmuOKAZl/xk6DrOmNGW0h7Gq9Uq57fDfi4wbxkZHKiCbRJr2HgYyrX3ljAm2ICYz5N0mcSa1CzgmYXzPKsjX0UBDNPBneBNvKiSHfLFys6tN5/nLiW9SGJcnsKQoR
dJALm99oJlbWIUAK7CpzmHqWeLXGpRHP3rxT5hii3rYaKDtxsgH65h1v2PbC9gBwLk4oTEX6+5UmixyVlQQDV8bwHkBoNjOFvJNR7mpFt207LukoofKOhWUsW2bfG5Wa
PAB2/kNlWR12cUMBTmPU1gI/QQsfNwCaeoNHp8y/lUMc2U9N0jymjkMvnGW9s0k00nfwrbwkfLUJ+KC2VuTnrpiHuaz0KTOzc4Pcu0+cneEluZCS6C3uGrvg0f4AvqQa
UDgVEGsYhYcXZxuZdnDz5K+u2Ajq72v7sLnJQfMhXsnOA4anbSQ8is3GwKsDyehsYlpeuco7gOk0utaPMGfgRcvyyQVIRFwOZxTJqeI4LuRBKOBsiH/t4d5lDp+EnUz7
e2+ZRdxYl6JUY9tCTd8l2JumJWieWC8ZJgZeirzAPMggNwI9/2ctd9YQRSRDO1YNI6RxHNwmt62zt4XXA0KVCpKf5o7mFjDEj22ZXsNJAIQ203gHGKD32JXG4q0CvP3w
ccfiOo8PBZjoWlcgdivzs1/jMtJq6kUo3++2KGZn7ZACe9VHkMpbTykH1QAzVcraFeHUs92Ludc/6LxKI31CxteVAMR867NPyhUStjIubk6BQeY8DuDnprg5tVMGRb2S
COWqRjbR/sRrxmNTuuQWexUrd4Rnl8wjOL9thY6XoKmG7z78osm5la5Tn3bVdX9YvnkPwr9oIgg9lb88ttsBi/ZSStt+ZK/cVUBmH1dpDlKUKyTfmwKhMQsWJaA48lz8
7Y4kGS3OIncg/FDI7oFze0jNWlsFcBD1xEOL9EszFtTU/msTv1u6SwE9Zpcmy59iztZEc7TPPDiwdSuABkGSHBiaUd6J6exjmyLQjEBsaazsHeA2LCZg8gzb7/Cs8+MD
O81NdLBDGVLlCIwEAKpVA55wHI8EYhLWUnZ1JhCQ/OWqAHOs1zKAntCVNEghawK1TL8ZE9AfGuHPekl20sALlzDYDo4Rf8wVRUtKI+qtQjrEi6KADQJ2w+QQNr87KRqb
Ns+VYRj0vJjm8rcE4ogFB7rtvKvPSsapHdwdMd4EpeUlXhlQF2H0yXRSNf9utSmwWKIz9Q9vwx4R442Tc3bJrwdJOaM79wM3Ik9yRCkidk9AY87GXh1zjNoa6I/aQNl7
Y6To9q0AnsdqfcVxvRJQsrPqzge+g22Bp+dJaQJvBsDz9+N1IQiYxFk+00ZOkx7JRnbv2attIpjNpKd49EGO6TbTeAcYoPfYlcbirQK8/fAfqw0r3dbowBu0dTQrk35b
OwrLUQIm8jVzma/03GBkDZV4+/Gc09NtZJWF5RQo+hj5ikFOhGAKKFpRVlGU1+2ZGDxUoZw/IhswLzA1zwNzLO/Ik1EGDfxjCGQZLO9fF1wjoysb7oyt5umlXqPn4Ipx
fXDCygJ5J7B7ZnnhoMsX8s1vChPqUwkIHkiEbE0r1jiJGueVKPori3bxXB3duJq4mqdMwR0MEKpM063cMUZhlfmVnaB8fqTw8xwRLZzWuseW0kHemAGFYeUh0nkKctOy
AVMl8gkM8yQQ3x5pp2uxHUcb7BmZaqNnC9JhAH1US1zit1dTn7ZnrvSZ7GRhjuozOswbmoQKQ9BdBp+aHwdJbTTZqMgYIgF6iAXYtvZYhnx5Iv53NGmg7tkz2U+gtjPN
8dpWiDrgzkocAn16j4z9/kIEm9Ya+TsJTV2yUmdvz6LX7YXoHlCeEKOzuHRW3z5oHEBUnLlS7LJ2FfFu0UR7urZCsKAXlBAp+8uEN8trv3GL7/tLHUPSEUkiHtDAVJd7
2avVza741t1OmCvxDyafFXBrTr9ZiHzg9PoTdeGbAdZ/KL0MmduSYwzribTPlTGrHTOMTfW98KCjn05UnIpWkFzzsg5NyAtJpOhm36VgeNSYraNMNTSbFazVbjUtK4id
QYsfZcpP4w05EJ4R1xFatSa8qayw7H1r43fSDmjLEah7zYH/ccU1DoEJMEKQv6lfTB49BkhaJEeitGtSyDxwdGJu4OJ43r/pgsYnaHd3zJJibuDieN6/6YLGJ2h3d8yS
3k4AMn7ry/1aIAuGfELsg1zzsg5NyAtJpOhm36VgeNQNPRKdgbR/ub6Mr9AIDgFw37rtGO+b3qq8hn5BEIEXHpGJbv4SjrBPWtjlq+SzwuK3wCJ6F99kzgu1qmXsny3o
DFbKoxd0vGchXuTzK1W7UgffUxeoJT+3uS1lOzqfguA7JsU+nmXh1t7+NZ7awQ53fBIC4YOnk3IONxLTw6osIgD+lAWm/FSUqjwO0tSswieMLBIQ9f+GwhZ+8sctuCSV
+umOCFv5PRFwInhZ4QtL7CQZTZBmNjp6khFiDG4HYnBhTjGaKn0D035J4RFbYYgMr3ZxUqCn1lLs3mxXuxfziEE2/lKbfjpBWzgl+CqtZHbuqnzEcQOjslY8W6gaoWJJ
MVPqEGhmyNq0LEh6mxxGk7TSc1XC9WMrGJj5qKysyYxmTj482Q+Xl+RRrdsSKTPsZ/9+/6fBU+roxKWahPD+QdjEvcpJHBLdnAZHPAEtVdp+EPjXVxV/1+bYjWRuBj83
kzh2vQqfu6Edovh2TGTlz2pMhgOicDReRo+LmgxpF/rIYNMHxg8q+r4nukrsIBBoXtz2fFacxULB5FejHsD+IXJw8Vj2iC04fHzP+xUom+mCODDmyYYU/ntE/T3k7kEH
ofd2J7hsoDXfx/tZpiaVpNp5b8976K5lZjA5YkBCsZ1IqxJHJ8D9bsiwrBfr7jUsVAaFBZVcPEm0uZYD3KsvsCQEBWPIddZyb+V/tOkwpL+LuFufTbE3YAgvC2EkfOmS
ZxRIxHGOFK5fTAtObU7zeViiM/UPb8MeEeONk3N2ya8VxXbHaM/eHh5B/25CWXlHwwGWb67cRBpzFzWhlUDTedv2yrZbIQCHY3y8nboRbUY1/pZyE7IDitTx/g0gE1RV
ENKrTdeZFCY4ahOSxjUWWcqIJtEmvYeBjKtfeWMCbYhnHXt0195sgpI/TPelBiBIjQKHvrz4b4NsndairJd5gzXLr8VAhPGvrXQys1A2zLLKiCbRJr2HgYyrX3ljAm2I
YqtMmuOKAZl/xk6DrOmNGWKrTJrjigGZf8ZOg6zpjRltIexqvVKue3w34uMG8ZGR8b0qqSjGDgcV77iDxmUsdMuva42DkVw9fAapLLIvv22YcvadVb+2/BwiuHMRDZYr
gbjx1FJxyyawsrVS85wLh40Ch768+G+DbJ3WoqyXeYNczJH/BEop9tCQelApxypD73YYIoCmPBD7ocBRjlBgsnA7TxoANRQLWoGxlHydiQemp5TzC+nmehOh+1arBzAH
bupnz73JmSSIv750IvIxGAZZL4JpkPNDCeBhZ4t19lw5KDifmVHWVEDeMHlvC7lZTQz5NocRQlk1KQwEjZx+4etXqsWfhXA322FvmKuU8Vfph9IYTEpA2xB6ygH3iTqJ
VFz5oI1uDUwJOUCxKo+IVfmiCZ5A0Y1IJz8CdWqwZyMUUu4kG/ToS+HpYPGCYJP+/OOEp8WHHy2CN1XELF0o5W7jedawT9EZ1i2zAJ0aZWQhuCZJdZgH4xGa9Jj3k+Qn
+Di1VzVxHjwJT9uAme0Q0EHnGrF2uYf0te7rqFAc0XLum9qwwmx4+rOPJcGJ/ERvirSuFShYByvQGU3iDr7Grn+7qtPnWC3WKFs5T8tQw1+9CvAkd528zOZMMX0xXIHM
wapJFD4lnaMwtld0cbJ8Z8s/ltSZEaGOsrnc4+Hu40zyHOSb9wD0dEvro7+oUcNOw4CggH4roKn1a64DeGbxcpHC+gC4+B0+/xiHphpIRhm7mFOqDifoUiObnYz+K1Wu
HlWzWHU8Cyje+P5aw5yje4z++dRTErPjK3GLYFlEFJPGAdOOAv+uaxmhd+lFdqVXQjmzwB8/PpbLCdfexu+tk32FEIO+GDxP3mLTT/YC9BtzbY8ij0ncDKJeQCUVrmyM
lTLVfViumUjtwbLygpeRCfda4+2Jjxac54CvlM0lYdAn3eb7Zh8N8z8FKFD76r7r4bTWUwHD4/XRz7UPajxg5WmTL/Bg2Ij01sla3w03Imkth3Rgu1DyNgIZcmDcyFC9
8nr1eBFl4ZLEsZ8C8jU8k+XXQxAk1s77SNCkcHY2fZiiLg4e7wsiEgfFpHEn2GgjTzjVkdD9ZusiD1yGFPKcRW91TJrjVUy3LVaEtLamovVohzpDbLM3otZJ/qXI5UjK
b3VMmuNVTLctVoS0tqai9VNJcmYsG0miUYsN1+Wx88KddI2SQlrfoHAGhUW/Qptt6KdsndLtbs6RxnoDseGp6AjLQgBZRpUT2N5WPYEj0614yBMEeqEZCCVjflXX5PKR
5w6ClIzX4b2SZ6VThR414GSAM/zm3q1IATzvCj6vkQdfdyFAvgItYTPjVJpvcdtS+idW6A6QYeDjviaI2VOM2y7W1t5rce851rRbPStrXMai220joald/NVPHVREGu38
FqRFModAxRnl6Ux4Y4ELo3C1d71rm4eq7XVouvgwZa7/mM3ruWK2/a/HYdRYhIL+UdP0vwS8crsz4FGGRZHt1xTLk6KhA1HjtW5IFGVlrLPjS4sAjKZ0SGXSRncJBfIi
jwR6bV55eDUKNGavjxhSCYHWbQUNG8GyyzqigTDgbfBwtXe9a5uHqu11aLr4MGWuRUO9i0C89bVCE15qKHrh2ONLiwCMpnRIZdJGdwkF8iImbyF1lQW2eGNW7ZtUnKXF
KxfM1+R8NCRCQorBqC/ApgNXqYoLeBu1b1L1YUJCAoqKGTTg12tJrIVCrT8VAvLpRJ1wT9RyrKSZkMcecsI6yMrSZw9naEvzqmJFt/gb2ZWQ7UC2qD3lKTe6uOu0/TfT
Ac4y5oRd5MJ1jTWPHV2WLVh5wsWuG/q33x4eOcqzXYG3Scxwr0u1nKw/zU3lIKU/40uLAIymdEhl0kZ3CQXyIlXuLz8v3xpkB8nh44voBChbL3rheMZoTLgkciLcGlOe
QX4u1MOpy/3olefrnAZ2HGdI1g/Dp8PKhXnHndE8ExjJhRQfEBS9Ppauf53qmEu3oYHebPJgkW5TrxedqRzZoqWjqlQOq+T4HLkd7feq18bKzYL1TCiHrTrsLP0Pebbn
k29ZIwUTTPhlUbS/HvJebeaLfEt98YzuZKcvZph/w/gdoATaMtzcQXhpNaSfGgkyPXcw0gFL+x0I8QAN2OIrD6gsJ7ppa5zdCBPf8YSbGFNc7fnFne8A5DN+Ry9/odcF
PXcw0gFL+x0I8QAN2OIrD94IsE3JAmSPVr7OnVtT9HkjT9bxrprRHz3hS0zA4G9A16wX/rkmWC+t9vNOlUgw2AHkuYZ265xXCb8hjpFQhilvYVuIFB4m8EYD/fWvI4o+
NxFlWzbmFY4875Fyskp3rHofSMbrq5Nsgr6nVccMbhEjT9bxrprRHz3hS0zA4G9Agqxu6dEZh4+g5vtQP7oicVFjXZWvmJ9GhibaWE9hpP2KZuVBTd5qHEFo5ZUAvt7y
Y+2V52tMw1+8IFuIAknorIZkLhhiIyECRer3ZfBw2M1afaYEwwu2vtthXHDvQ3HGDlg8wAsTwgsiPZvrtOKu9wVjovR8B7ut9XF9+kQBKvjbDXvn3p/izVCOmJbunRM3
ZRru3MdZATchFyItRtCgf0z2E3GnpdLHBn5ZwaoNfbUVK3eEZ5fMIzi/bYWOl6Cp3HhCXqFrVRrLEqNT1d18pY1dmbJTdn5xFqDltKKOBK4fZ2+JXso8fkrkF34Tsjtt
kpFEAHvAxIcZJQskbG/0VvjVQ/TvOtPKLUr4unLYIyUzHap0xxKEuXnGGbb4+9q95fOgLGHbU1L5EPpjgggvSM4PcvKgxuEMi//qvRpGuxG49s2ZGaZvLyE4CzSEwP6C
jOh84z0hyVVQgF9xEdD/stpF5g6+kBABAL2rZHl+5rp9Jq67nZCoaKAeIOa5kZU8Mx2qdMcShLl5xhm2+PvavUV/qG05OnTwqYSXV87NezppXG4c3A+C0wt1bw7esD9I
wpx2ujZXFZHzdkPruJJLlWxs+i832qEpfMdtKL4QQM9VHNEwjuO3tUV6m7vRGUtyBTJcHYjhd6fKG1j3nHDzNZezNjj0XmKI7f/5+BLp6loMFWawRfvHc70B3o01CvwC
uzqrcPwr4d3hCpRC17g+UX072xVOYgICQjgqyzKjXgUfPglAHcCqd4tFGZSh5+UFFC39lISk2EF/V6bsZgogXXFfNVC42VzKhxt9zjVumJQ9H2mZiOJ+k/h2P2pO/r4P
X3kxbjITxoyYzoAgquV2G3bPjksFwtRvKHzt4O4EHZauG01CNsNGqgRbQ/V3iHzEora2FFctOE8UK3wjobCN6QJW2AJKxkzQkJBOGlfO3/YzMAZ5aut6BrFRHpnrdA15
FSt3hGeXzCM4v22FjpegqUp3I5Vi3fnnn8u7lINYw3zzqfuXfGBYbUo0KAXi+m8f4AMMVSAJDPx3wL8stvRAWstYzyFJns3fQ2XvGOZumkg0donda2wIrJHSVoTyef5Z
ytJnD2doS/OqYkW3+BvZlVs5Ii8hdReIMEo7+PHPfbxzHivAqKL5sx+0xNkvAPANy1jPIUmezd9DZe8Y5m6aSOhMtqi7hrGpZX1tjNdeVdFW8DqghSiPwaRKdGR8cXXF
RX+obTk6dPCphJdXzs17Og6PbNBdrRy+EQRR9YU4cjU96sNQEddbdKGX73b7Wb/ZoIezdO7bAS8U0Ygw374tMxwjD8XZqNT5w8i0cJfBOmSA8qshhN0tNpxESGapGjW3
ZRru3MdZATchFyItRtCgf8ksAnQUbelvvfOVNTBE2wmztCuflcFq9LUPtBier2SwLj8ay6Osz6I0b/dm2f5Tk/Az6K5bD+bZ/OFriefwynCFToT3iDuY3L5pxzKgMi71
0aoTaEookCHRgQBzTurw2j30iD4F8TbgxwFYP57ADyqbDd7OtvuK/2/Yu9cjNEosJg1ibuSGn8sg06bdksahKTNM/Pfwe17gc3bHlSZrxMoiDz0kCWRwYpA7wim2sk+8
vvjpS4hZdn77vjGpHqhia8DwMv6P5N/C4egH9gSNxA3zqfuXfGBYbUo0KAXi+m8fdxe9pO02pFvOckGxFLkqpRUrd4Rnl8wjOL9thY6XoKkRODiaI5iIQDGNOP2p1yuj
Q5dKgADt2M+RhFeFnR07pCswi/netMNTr2sOVjrXJJkEtQc2RsBdDVz6ZLHyUxdlZRru3MdZATchFyItRtCgfxDtEGBCvXA+gd6nDVFLnD7z5HSrtbg6gOfBSLxlfgqq
dB2OuGVtZxM6Foyw1GBd8rkCm8tBvOQca9LMMHOhr8kN94iTC1tlfuSUHlVV1wiTuQKby0G85Bxr0swwc6GvyYhCyuOxELLAZ8bSNin7WFd5Pb/JSXo4V0xDwPdMnEsh
w1suIcYf5o9w+RSHMNJp1f1ZN541VLM0Xv0vZej6MHcOvqx973XjfBXe0Z/H1pvXS1PGBZoQpKCbP4afa83N/Vh5wsWuG/q33x4eOcqzXYEkRcgoKW0GbOYSpKpar/j2
Ep7/rpzJCPNPHtdfrlp9DD0faZmI4n6T+HY/ak7+vg9l9AMnUCTG6xYA6RJRivpH/0hZQfFjIvB7LH/yzdYDLAVjovR8B7ut9XF9+kQBKvhTXjSrqfx9W1ZIxVRvBc8P
Mvkd3XE+76NAukNXzey9mWfXRcQT+IUXYk2Z8SYeaBdwtXe9a5uHqu11aLr4MGWu5fOgLGHbU1L5EPpjgggvSEtTxgWaEKSgmz+Gn2vNzf1YecLFrhv6t98eHjnKs12B
IXZablWFi5GlUqK/wVdZaWps5F3r4/eOJ5IYPdA+DH/Hp8wWnDAjcfvhPrQXyulXIyEk4bQ3WLN+w+TBTdHfh75m9ZWnQ73MhKuGubdNwdAEHUikC/Ixlt8sgJ7gJmLa
YSkZof4QW9deM7MDj6Lidg33iJMLW2V+5JQeVVXXCJPuv8wdDMWDsStRJ8uAeuzmJbmQkugt7hq74NH+AL6kGiMhJOG0N1izfsPkwU3R34fFSvzN+h+6tEuvTcDDdDQh
Lp1eTstbA7M5Hn+OiHsCA1h5wsWuG/q33x4eOcqzXYEI+iUiGgGYjHoeLgFf+QRB138JmrxVKRKGUH2AsswEumcde3TX3myCkj9M96UGIEiNAoe+vPhvg2yd1qKsl3mD
Dw63ngmEXdWgRI8hy54Bo/y3eSEDSf6G66H68kXVJ3RAxWS0dU5XSPGm+rWQsSmKm7OUpyqr9qjffPe27Ox6AsfN2tp5HcfmbKEzcwXh6O9wa06/WYh84PT6E3XhmwHW
AcTvF8gwooMKmKArv5m08N5wXG4D6ychaICUULjxIn6z6s4HvoNtgafnSWkCbwbAcVNL5uoVyWOyfzy+WoPcz0siLt+a8sSjtJu43cym9C53gK4/wChqFliJXGHIobED
2/bKtlshAIdjfLyduhFtRvNsOBGl+w30PbDnxp3j+4rjhCzlLVyoTWIpRcyixMElivOe4/l8ZFWmyFZJTJtcDWJu4OJ43r/pgsYnaHd3zJJnZoA12sIVcFBBJq4HZ8d9
SyIu35ryxKO0m7jdzKb0LsnnwFUeV+nIj0ZSulZAMGdycPFY9ogtOHx8z/sVKJvpaEBAYmrE4d/1aOxlVlIQEaqBSMbRCzcxPOSvjyeIN7XDfebUsBFoQkaV/7M3VcOM
zwFoJdrzm/GGwvRO85CvPArjSGBk8bYz1G/l4lMSQFsFJ2dz/UzDkUVplcBdoNPj3TGnbIj9fSpgS1yM9aYKiic4CUzJ1tcVZcw7bBhoaeA/9XMcOAE5Leb45XZt9Km7
DXhyHYDJlJY2T8b0jTqPxZ81THHxO1IqHElkWO3vNkKnMJP3w4u9FBMD4k9x/6a1wuFbpNeaeJKP66nqS66CmLlJn++I2nr34CUDxN/37bvXfwmavFUpEoZQfYCyzAS6
UJY6uWUkEk7UQimZGt+oz2vpvYmi5QbJ+AzB6b1tv22rSh8vVw4zdyiGQyU1lt5GQbACccEll1A7qAjmWM8Hsz95jirKO0LpkVA7xeeAxcCeqeJ6fWFRA+GxKxSB1Hw5
Ia9P4jfZtMWcLInbxEO6pBvBQLHAy6x2DzkQyM0G4mA4DTG6mr87zLygUnF0fTXdrGJ6aQdmhzORWUc9Eu54pm6Y82hWBRuhQobCYN9ttZrRq7Y6eGwp8qmrJDWGhQ7d
K3DLtnBVvA1gjXBRM0SI7gmbzPExbhQpAgTRi/SqjyCO9kkm9e/xyOYYU30bMI75EMvQ7cuUTt8YjOG4X6XSpjbTeAcYoPfYlcbirQK8/fAVKIeyQoKUldb0vmH1luWc
duRERHTC1rah4BoDk25mRxpewWXWB/E7qZRAuk0ixh+rwXGpZUJuCLu+B7XrJgx6tKoVvj2KnHpU+8Cf66MEIVdftnP0vfzSGYHLXCezSPPCFE3pOmNnshjsgP2fEB16
i4gFkc6+uR/wRaat2KqdUr0OAht2J4sJW6pPArsCeZmxYfXqIxjo3NseiQFDSst5HL75EhoHB5eW5vXYt9vzDItlG5Ew0kEi1HUSNFn6amTXDPzOW9Ys2H6KS3GRHAMt
Ej4mP0dP++gi0j8WWccgYilNuoUWukNb8jrMSESijVfcpxjbTtEsgRBP5Z2W558Cjr6vTM2aVfipelRHffmQhnfYWCgbHJvTI7vdvtpPnMrK5Nx69gOAhqsX0zGgP1Sy
zQWyTxkf3I5h0Myr4u88veSDR/bzZ+/Po0PurHP2mnde3PZ8VpzFQsHkV6MewP4hcnDxWPaILTh8fM/7FSib6SGi1tb8HsKmhl21fXmKh5WqgUjG0Qs3MTzkr48niDe1
w33m1LARaEJGlf+zN1XDjF/LaQH2Od4954mrqTk+iRqDkIYepfWOjDJhRUhhLj5pRFLZcUMOqu1bP7hiQSiRXo44mqhmo/bli3oNE21FLOHw3Vo/GZ6/DKZ0NKV/Ae9Q
LIGmqlX8ehcCqqeFOYiQmrJKLXwq7QkZCEOQNFsN1Ne60UH88ZLSHFZokl4sBXX2Y+8XzRuL0QGDmVbPwo7qGo+pLDh1aa+HWy9b/aHr8cHt6tLqEEl58l5f8VU6Qlsp
eugZ2+pDPXYw4zX10IfVVy0xpyK2xm8D/LDceBUsfc7Lrt+ZYzJEeEemyEsn/5sIUjpU3OoSC371GAWNiLvG9itpx5K52wV3i+CjixQqcyIAcmBid61FsUikVpKpE1wa
MM06zAsD2tJ1Gn4dkASwNgNPwuokwszRetD34YKLoj3tBfD1cNhsA7nSuRhZSPBiqAxg3HSCIwFtCwdHVSs5Rf6rA3cHMP3pDAibLLfsgGRJo1tiEzoRxqJ3BuawdKdY
REUW0A/ECTT0choTBX8KXJMzy/SQM3WezP4MQqIxAjxiWl65yjuA6TS61o8wZ+BFeeOydXEwpOEsxnEMq7BU7LFzdmAWJin2+D1WKNfVn4QWo3IS5dFVuBrypx2GbVeC
3xDTjIFfQfiTuF1UvJRAuxZt54UUrnNreFmC0OrmLuYDLEFtmdnKmnjtcvRt8KYQjXBJUItitJSkFIibzpYm+dZ2PS8H36DETzePr5Q/YLkamnW3/x4T2hmCTlSFI3qc
k9eFxoGmQMOV/U0RCNKn+BPxYDyeQhfaIXqmCkci3cJWG7mfgYGWd3nuKw1OUxy3jQzPUXgfYuDIqT1NsezZvqFMUxusRTDfS1+ZjuvcqmB600Zt89Fym0TmdFLAFqez
JryprLDsfWvjd9IOaMsRqIVfvllyokCNmZAjnZREe5Vcrksj5ZKt25sSZcv7zCStL00+VoF00p1m4QPt4caPxnjJJ4OpZvEx50Dj/WVRFpmtV0c00tY+HWUU1Ol6JQWK
+TxSxhbkps3ar8f2leecWKHY9tQg6QKbR/2iRrFOXnBu4XFa0c1Gzb4Q11NQNUZ4mazGpNqFvIb8wzDpz2rQIKBNjNOyLokHwB7jXbRsCvgtyCnIpXh8Ww041tJFbUI4
BQLZ7Vww8Bx4MHrImwE1LM8T9jEA6Gd7yeJozKeUI5pMc/I05FaYudweIBgw8UwvuzAwDsOn2h6ucH8/0CYWPNOZrTjTXjjj+CPAU9cPFuwwHaRUJPWBA0rqkzAnZnES
4kpNnTsHIOKa8hiutIyBa9TekJdtfpkfWaS+1bbGpchg52PIM5QL6qHD5K+cx7Qf2m46tnCc5/9i0GPK39FrB8GJl242KNDCKcUQBNV1jX6FT9fB8eSjznfsSg00KVC2
Vhu5n4GBlnd57isNTlMctxVCN3TcMnXKa03png3KsPlULyUaQccD0+1fvCyNEB/ydHZWV2hdxX8W4OKc5HXgPGcde3TX3myCkj9M96UGIEhmuVFFDOipQ0wMwJTO/MIR
2KyLNew+iRKoyhz7g+PQt3l6yzhVLlcXtxiohkB0h/Nm7DHf28NyI8i/b5iyxj0e+Waoh2CfTvEXRcGyNkvpppBT1Mvb7MB2H0SjRNMNyL3zbDgRpfsN9D2w58ad4/uK
K5oFaeiqv1eeCf+/ruV8Yl+BM4f1ho7a5UFmfYczr8tN31NwfuplLS5k18eIh3MZP5Q3wQq8h+L7os3AL+5lg3to3MFSbnzkK4O2D6F98Do5rgVRMkuQJ4UV5axzFHOY
jeI+mGtiXR+J1a1WMrPTYSSNhsneWrjn6ocLnmeTYp95ess4VS5XF7cYqIZAdIfzEJuihxIoZdIX7WIyl9c/rrZWUAcqTWJPUg4Pj3Fu/sjiI816gMcPUBeoNYpCqCU1
VvYI7+QAxTLIyJ5ytC15EemjMgrFmrJCEL076GISCIos7CmM9E8s5GWoQoeMl8YtfLsOX47/byY8lDHFS+LQXEsfiexKfOWr8vk7o479HVYSJFgvomH8TwNgovjC+jK9
UbwAsmNfPYVBn3c/x4wCjmkTpKEwP89YclJ7sYGHi1qj0NpHB961hhHzSHPnU7Q6866d6Qw/1GyShElsCQmxIL7s6viGBtR8fA2G7rly7SVR8v3EIZj9cxlNMVndP3wG
beBwki9HpTvP+jb7UK6nD5szsX6G8KbWqZsktSg3k8IButiDTzz2SpGjn930fmK6ntmo/7oJwbEl4VqGri3sKgQ8mGyLag3m8rPXPnlg7agFVV/hDeUtU6n67HkPhRvU
DANv7qIf0Cqi7CW25RXqunhRWBBzrmYuy+mv7t7zxs28mciiATaiV2lxR92Mf3BrV0uLnaJlkZv96SPjDychzR3Qp60fFs9uOjurshYVG9paSC8YyBC+sSYYuVh/Qo4n
vc3vONugujbqXQFTpi4XMrUSRl7YmxOjAFZJ1Tw12HXjXdvSwKsPwaymJYaUpJqL8v0Ih9rKzwNgZ0947id+vnhRWBBzrmYuy+mv7t7zxs3MJd267ttv5SDhWcS0S06e
n4BTEd0JvvXCXHvctoRgKLyTykqI/DP10c/jR68exxNZpnqbUKp1doWl1qjUOSbNU1V1n2YjMjUGUV1cVMyEm66Fi7rWaygFF9mW5qWSbKRMtEJyUNCWX3mLenmZOWE2
T2Zm4EYcbM76JNH/7w5zu3l6yzhVLlcXtxiohkB0h/NxWnIYRPMNulq+evCIzuo78WGpcAZ1HammM1MB9eeNc/sEhiT+CQsyLt6VABC98I5wCCsGscX6uY69uODSBDBp
xONzOoQU3YuJmggeWyKEQrW+SnaiepOjejiJ5bvbY2GG+s5mfc0Okp0hWcZL1pkJ+RJGbCNiEhyefW5F56kI9JCXpA7tImgxVyRo7p1WJ1gnz48UcfAUDy8m5MjqICl9
beBwki9HpTvP+jb7UK6nDzxePqAzYE8H0KPF8XARKGoVGYgLzKndlb9Uc5SNcLwAyjx9yJ3ZHx1GIAF3DanAj/kSRmwjYhIcnn1uReepCPSQl6QO7SJoMVckaO6dVidY
B10zZ76DizE56ppmrRmOyW3gcJIvR6U7z/o2+1Cupw8ZHQM/M/JZDf+hU7Drq4q1L8t1RPxJw3m163vMAtyVXwdJOaM79wM3Ik9yRCkidk/QYPgN4h5ZUXRYOWvks0Nv
pa58sJPAu/P2mu1LKXldRB8+CUAdwKp3i0UZlKHn5QVuq64ERrR/oItcEjuZq1MFZ5R1kyxoacl67r8VlnFmX7746UuIWXZ++74xqR6oYms8w6jq3wOTZMa4vsKf8Aey
t6CbuahMo7ZiIYMZJ2ocTHKQDAVLaNwIcK34oRo3h6+kU6INqtNgQeas/q9Jh2oLtG4Ky8Jo1VAwqfpk61ify//BkVvHrHYYzvCxn0uAMdWkBR6MrbqsieYWviDOinCL
Ix9rpY0GIiXSkUp77XzVZqHY9tQg6QKbR/2iRrFOXnBaZUA1qBqktcIgpYFnpQbMlb29BlB/YJWQta/18HYgj9aKa+6wcNvIxDjX51kkaJqtt8F8DIJkMFl1VuKlLAjz
d5U30bhGeMtvIjwFs7c5vLPqzge+g22Bp+dJaQJvBsC1JhqwMj5vXZYYHNy1F3ag4tfYfaZei1zguvys+5NVB0YsS5cQO3Dq4ERL4T0DtpAmvKmssOx9a+N30g5oyxGo
CacpXmM9n0LwzzIAjMHX/F2HCq+G+XPF0NlH7Y76LjYcu09gZlZiPM0NVkhATLxlodj21CDpAptH/aJGsU5ecAqWt+8Qyqij6AGDesAQrTV4UVgQc65mLsvpr+7e88bN
Hdq1XlMN+ClWf6+2niW99fm4hrz0hOvokY95V53GBgx27zO7sqVMZ69RaD+ZcYqUGvsTOm52p3LO5axkTbFnnQIrGWBQbDVs4Wu990mfQ0k/GrLc0x+k3IvTyDwoeGfZ
GvzgsAuMOzwMO6d+L2CZdqHY9tQg6QKbR/2iRrFOXnCr53ofO0fGaTc2hlYIzJ0dqjJqYyDySnealSXY4HKV/lYbuZ+BgZZ3ee4rDU5THLeaZa0Warz8Fol0Pbs9hC6M
eXrLOFUuVxe3GKiGQHSH85TPSxQ5OV3pn3j0I3adBYgCKxlgUGw1bOFrvfdJn0NJKsEthaLjbAOaR+4hnOmuV7+hr9rMBt/YJtTLHWoQ3Rp1siXEpye7BR39rSreNMDV
RsAFiAbC6hvngJAZ4UFnEKoyamMg8kp3mpUl2OBylf5WG7mfgYGWd3nuKw1OUxy3mmWtFmq8/BaJdD27PYQujJUoVoCc0FG5zuY9it+Z9piUz0sUOTld6Z949CN2nQWI
yhI6ph5OKxCFg0Q1pDc+RoEIU6G7yBNiKx/361UO/MdHRQKQuarnyUa+UCUEjAv+1opr7rBw28jEONfnWSRomgjZFcvcb4GQblcOhpX9fw2fga3z7xftXZFhIhDd7Yhn
L00+VoF00p1m4QPt4caPxnjJJ4OpZvEx50Dj/WVRFpl1jDvbEyZ/b3r9mrG40iGKYm7g4njev+mCxidod3fMkqSLf5Ic0qtpnTJlpjl42uLugw7rF7wkt9IRl4/bvovq
0OGI2xjlckJjBsuYUPHZTHWyJcSnJ7sFHf2tKt40wNVGwAWIBsLqG+eAkBnhQWcQLvE+KEH5/5oRoYOGepVAHg+N327w3X3Gj04PhMjF0UrAKy4DI0yQhrmao7lNbVPx
ZNLJzxEWQxSFqJEcCcWWtnfqGyt7YqtpMq6HCNINOg2F6HLZ0smTUbbd017inmdaL00+VoF00p1m4QPt4caPxnjJJ4OpZvEx50Dj/WVRFpnY9uZ6ovT8Qa3gtVULR3X5
/zowf9w+JeqKUpBd08q8IQkwI+xns9JBXH/rkbTOJSohXw6uXly53PjolaRI0D/ymM4S4GP0fnbtxW+M6dM2upY5ym1Oc26G/IKUcihl67pfxD2QS7EmhakcnXZAOxCH
ab6kHh8mwoFBrcIBQ3mFrrPqzge+g22Bp+dJaQJvBsDtUG/7xQDY/16q8vG1O5T9X8Q9kEuxJoWpHJ12QDsQhydfsvbkVCQTquaoHH7VPGi+RS293MpOkXba9mKzk8Iu
ll6aGa3StrIGnRgXTAWSD0BAhEgWSiCGmbGEevVOmWmaLLfIBAaUMawP2diJcKLbIV8Orl5cudz46JWkSNA/8pjOEuBj9H527cVvjOnTNrqWOcptTnNuhvyClHIoZeu6
X8Q9kEuxJoWpHJ12QDsQhy3IKcileHxbDTjW0kVtQjiz6s4HvoNtgafnSWkCbwbAc+xyzdd1fngQvKscIT8ENNvNJ0t4VgWQnTsDTDujSwUkNQgBwMr8BLZ0n1LSNkRm
cwUfQGdNDpf7xB7zxU6lsgNlO5XlOr/Q7eX4glp0QixXfU3DausIxILYlQpuW5ss5WUROPrvRUBLurE7fzIebcBzxhzS8JMs3NfZXrwD//QRZ/5zz0Dnt+XYeEgc1lAs
VB8e2K9tb3XyNaGbGWJCCe7Be/RuOYIY3CsgEOPg7JLgWnpYmjvhqGRfURB7RbLMJryprLDsfWvjd9IOaMsRqNmTCue+BgxzDFyMJ3K1m7DhFXmAbR6Le3mBWzt5QYgB
Zx17dNfebIKSP0z3pQYgSGa5UUUM6KlDTAzAlM78whGUoiIzlBl1elXsVW+2TcKUeXrLOFUuVxe3GKiGQHSH85TPSxQ5OV3pn3j0I3adBYg858TWybR9kvGeF42lTG4v
VB8e2K9tb3XyNaGbGWJCCV0NYEBxmgE68mkLpSPMlpV1aKjbnjNwph+4oy08w81THLtPYGZWYjzNDVZIQEy8ZX/vYJQMm0Fuzb+cy6CHDx3gfvDPIL44o4Fd03QNnc2b
N2Q36AzRQ8/7Y9/fcvaOo50bvupPSkv/bkE9dD0OoHJTtio4OVdY/FheevjSNUBx4tfYfaZei1zguvys+5NVB8OaVnaC1KpRI5IEXK/9gw14IU+NIMx6ywyK2jWU8Wys
+El9dNPTuBdFtAoOfPK/Fj7r3u+si68k31O/SMWrv+ITczNQi2q2jlYoXRAYdNWipC2WC+rken9jA5fw0Tn6eSy52HsQox0kGxppjLmKsY6YzhLgY/R+du3Fb4zp0za6
uiCm8njov2PnOxd1ZF1/w/ypkMsXrn0tRvqcYLOoWKT8CvFL9nXrqXZvAioIb0/7JryprLDsfWvjd9IOaMsRqBFQACeDPEUSlfQ+3xEi/0ihuOwV5Iuy1m8QbFhV4wBx
82w4EaX7DfQ9sOfGneP7iugttP+vWFtp8eBhhwp3ImvYoHHiI4uh3gd+N0ONAkmWnRu+6k9KS/9uQT10PQ6gclO2Kjg5V1j8WF56+NI1QHHi19h9pl6LXOC6/Kz7k1UH
w5pWdoLUqlEjkgRcr/2DDXghT40gzHrLDIraNZTxbKz4SX1009O4F0W0Cg588r8WPuve76yLryTfU79Ixau/4hNzM1CLaraOVihdEBh01aKkLZYL6uR6f2MDl/DROfp5
vmGdEs1He8z/OmzpvQFKInjJJ4OpZvEx50Dj/WVRFpn6UE8+C6JNJ0ObUAWb/RiXqVn5khXzAhvdHUwF9WLOUdJH7iemvQOlugNy0L30h2sgktsM8amgXthSy3oT1f+o
qOTzsHQk5is0PDC7KFhWI3q2jHqek+fokHjWWPSjMrvSw2UxGDfZZ0itArQ57R/Fe2+ZRdxYl6JUY9tCTd8l2PaeYMyWR19nt/1HEY5EHNqpWfmSFfMCG90dTAX1Ys5R
0kfuJ6a9A6W6A3LQvfSHayCS2wzxqaBe2FLLehPV/6hcq58TXhgCp9wo79XorcscqPHGk4W6Ro66f2JPyKavO2pT9DZuT5jD3V4HCyzzUxCJ9XtFdoHrWMocQkj5X3l0
UwCu+p92PU4zW7g67Aum+pZ3iowTGXVvbdTg2NUYy8vyVYUHw7lccA9EweHmI2TEeI4jUtPLbVAaNt6W8K0zW2DnY8gzlAvqocPkr5zHtB/abjq2cJzn/2LQY8rf0WsH
wYmXbjYo0MIpxRAE1XWNfoVP18Hx5KPOd+xKDTQpULYBxO8XyDCigwqYoCu/mbTwcRe2iVdpK/VqUzVBaAVpqEP2vW6fDFaZvDkhklymXAzAf/DOs1Mn02Qlwqo6oLhJ
05mtONNeOOP4I8BT1w8W7DAdpFQk9YEDSuqTMCdmcRLiSk2dOwcg4pryGK60jIFrVwpV/2rd4cUR38iDwHHKz/etSo46JNIh2FMgyDkdWK7WBmr7mOv2uWwAsdMZ9OgQ
xUr8zfofurRLr03Aw3Q0IWGDC8akFg2gqAWwaWrUuz1g52PIM5QL6qHD5K+cx7Qf2m46tnCc5/9i0GPK39FrB8GJl242KNDCKcUQBNV1jX6yKRGtE86Or3o73VsibHXC
MB2kVCT1gQNK6pMwJ2ZxEuJKTZ07ByDimvIYrrSMgWv4GO5ZPK0dT+zEgIb86x5gJW9VEdLhdlG5zR765olwsGTSyc8RFkMUhaiRHAnFlrb3EJAANx4/RKuM5XnFs7Rh
lb29BlB/YJWQta/18HYgj9aKa+6wcNvIxDjX51kkaJrkBJcTd/nSwByj5QQbHG/x156cp45rxA9jcXr/+2fTtOR1cTXrYLnN+0x6oQb5PiCHCiJaW84xcUjFkm/0tp39
+biGvPSE6+iRj3lXncYGDOXTnk8Gk47eP/vru2/KSdn8CvFL9nXrqXZvAioIb0/7JryprLDsfWvjd9IOaMsRqBFQACeDPEUSlfQ+3xEi/0iAl0MS7xVjCqcc8hq0NFyA
GdC30oHJVEbSL7chcEC7vqcF9pzbRTAWzUQ8xI3q+lKitrYUVy04TxQrfCOhsI3pAlbYAkrGTNCQkE4aV87f9lzzsg5NyAtJpOhm36VgeNRm7DHf28NyI8i/b5iyxj0e
1GBcgcK+SBbYRTFhu8BbtSgZQf5rhE/g4X5x6Kz8e/pIXjDN4gPqCIxW7OtyxgvrZrlRRQzoqUNMDMCUzvzCERDXuS+jCGv3h7oenQ26TX16tox6npPn6JB41lj0ozK7
Ix9rpY0GIiXSkUp77XzVZqHY9tQg6QKbR/2iRrFOXnDO+w3aKAsJGl+HCx3DWQnhIXKWAhhZ/J+dMXj5DEf6OajxxpOFukaOun9iT8imrztqU/Q2bk+Yw91eBwss81MQ
LnoQU1izhW9vmCcKlvo+1cy13KeJwLIbOoWXS6NmoT317u3M6qcndbDKB2J6xg9PoFUiSXKgmTqgsgY1JynXNKlZ+ZIV8wIb3R1MBfVizlHj44rRRXWmXeSLtTXGkr4t
JINlsVNuJB/69+e/tLPSfOPjitFFdaZd5Iu1NcaSvi2JTe+U0xiAQ4U/7vP+jxz9YPCf4GFs595XwvKx+Srzs4pF3VgqZXG128SEw1ZmpPNN31NwfuplLS5k18eIh3MZ
qRznql5NCBeJD9xVPk/tpQbm6UlUst71sXuC65pyJYI5rgVRMkuQJ4UV5axzFHOYjeI+mGtiXR+J1a1WMrPTYfWcpMOkZ9FMsqlVshjR35akLZYL6uR6f2MDl/DROfp5
dlsWm+1BnXjjbxLLwDpwClzzsg5NyAtJpOhm36VgeNQYLRKC1B6JVCoDVYvIFLu0CUG5/uvuTyW/jziajhHRynMGTn41CxKZ23uT6FdVu6yDklndUpEmPbcQaSNwovuA
R4O4fhADK4/Oc3JPkiqbPLxe/GfTMEpUbJtFwYKZxbLVY5LSjRTE0VUwi0575SOoaIAT+6h2/ykPNL9POFEc6vwK8Uv2deupdm8CKghvT/toY9EPHP3TP8Dzyshya/i6
i/ldmmH0JWpO3FUJeWzOY3KfQQHtbWd6JzZFTulSkltoY9EPHP3TP8Dzyshya/i68IziSWPVGXfDUC1f/J+IB0eDuH4QAyuPznNyT5IqmzyYjaXKsgkk9WoBbj7C3DjF
pFVecl86LywKOVxx6m0GGuocQSgc28wTmVZvVCcsfYSp+H/gVziWCJfW3Z05BRsLINOFQcclWGsDbTRDdk6WO7WMk+hs3ad4UDD7NbSnGdl0C50vbLIbbcfsZ8ae+9Us
aW0MZ4Qdrl2vqEExw5wscHQLnS9sshttx+xnxp771SxJYEV5wBZLzjmc2kibdNri7Nqasinvv7Wqm/PXayWpb1jhlmM6D7YS/L0HzbwrMZls0IB2+kUxHojl05lKmamL
Cy+AcKLPRKgVqZnXr8umGg2xzZhnaa6onO5zrLlSbwo69j/L+juuSVXjPd0T9KgLwvgJJ7ZXPeNACHGIZ5ucLPHd1vuaWwz05ozNYBgDLLR/NzSZvS+dvULgKVgM07Ep
cLV3vWubh6rtdWi6+DBlrrGJZRW/P7GlZEiK1c8HzjOoUVvoEmK53L2KJIHPpDstFSt3hGeXzCM4v22FjpegqfVzO9rb7UR49j18ZAdK5jY712WCVXDEUzcr3vJN/M3r
g7V/SY3UW2i0hYydn43bVaXl0UNAFO0yZl7MyFhHAJFyWrytrD8FUVPSct1AS/0jbymzngLMW6igjn+CMznec4j+41bml+OhWPwdisz+wZpVm9QFYz0hJLvSVPqBA5zE
uH0r/smvfaC9HDXzW0y0FmG6ZyvPbBLkB7FdpSj08vo9Scqta6jxnDOsP08zfcMK84G6yxwNscMQ7v7Q0eIP1IR0kbPeQHVTgE8feqlLdLq8n3igUvTgJq9rvcScR00O
8kXnzNM6KFGuiE0KM4Ey7OBaeliaO+GoZF9REHtFssyrrJrkcvtFkJFGgG511EIKAlbYAkrGTNCQkE4aV87f9lzzsg5NyAtJpOhm36VgeNRxWnIYRPMNulq+evCIzuo7
8WGpcAZ1HammM1MB9eeNc/sEhiT+CQsyLt6VABC98I7AUyn0iIoktVGfdkXmTScx1gnlQ9vkKsNBFsP5W3pFPGskNRFMx5AWhdn9N5xx3ExPLfobdspQgYSKIREv30fK
ly3QTZvoamLYR49HRvpPmsVK/M36H7q0S69NwMN0NCHG5fhJxL1RattJPsgd1wq9Bp6n/WvKF0PK9Iga995+mzvXZYJVcMRTNyve8k38zeuDtX9JjdRbaLSFjJ2fjdtV
peXRQ0AU7TJmXszIWEcAkQEYhzxgW5yDN9C8hiCNKfiymsv0Alar2YzqSwjt/qH21SmXW52x0rxAa6u6iIeYu6Dpy6MG7zgSdwA8qKnfyrVsMriN0fXFP/FJeOjbTcM6
nSSqVw8/wHqSonyLA9/sWODibBAiDJuN8dsTqRLtpBPPbspkrCTwkoQcrEC0frXS/ArxS/Z166l2bwIqCG9P+8I0y76qbW2hzgUwo0a2FHyDSFvRerNEQpWpZKjoOAKq
fJFGx/kiBdBtky9eK5o0kRBA8YkWHGoy+WeBsLKzOWq4fSv+ya99oL0cNfNbTLQWYbpnK89sEuQHsV2lKPTy+ljgZSlBqtG+gycpJ/I4lIsnMOcD3UVl5U1ucxXFwY9i
M0z89/B7XuBzdseVJmvEypDHHxUoiPfHd43iwTTQUZCaldS9bTTK3f7HX96zq4Vdfw7L3OlJXtAeZBNwTotiUmFUIgay7Wrn/kYlVNX4qZ6ORwen15l47gBfpxVN0LuI
tPdIaG3kVHM0t50lrCrtPswl3bru22/lIOFZxLRLTp6fgFMR3Qm+9cJce9y2hGAo7j7aQZ9J0OcK7Qj79ZKoOBcgMktNBrfZx+7ff0TxBrBKXcpqdW9metrhxY+1aLZZ
amzkXevj944nkhg90D4Mf89uymSsJPCShBysQLR+tdL8CvFL9nXrqXZvAioIb0/7wjTLvqptbaHOBTCjRrYUfINIW9F6s0RClalkqOg4Aqp8kUbH+SIF0G2TL14rmjSR
k+dANzVrGPmgAV+a9wk9T9YJ5UPb5CrDQRbD+Vt6RTxrJDURTMeQFoXZ/TeccdxMTC5PduNHw6G+cF86c3KpoAhOtfMeUFnHlBj3ctnWwk3FSvzN+h+6tEuvTcDDdDQh
xuX4ScS9UWrbST7IHdcKvQaep/1ryhdDyvSIGvfefps712WCVXDEUzcr3vJN/M3rg7V/SY3UW2i0hYydn43bVaXl0UNAFO0yZl7MyFhHAJFMsn4tRXBuV+GAFxabcMI6
2qJRELsSM6nwPNhuK8tHqfMv0wYZBDkWmHiiIuRfT3KTo8NlBiQjMkN0IrB/0odzrDCutQr4IPdJScvIwlUBQ7qZcvRo3DYXsF9Lipf58ydc87IOTcgLSaToZt+lYHjU
TPgu070M8t7i2mW5jd0IFgK2ghuqzolbqNFwABNwTB6k5MnZjnxwDkv7h7Rj70GXvdcApQMQCV5NKfigNNkpgH9V5lnijLjFn4O8rkIRQ2TMtN+D7R+25UEuNrQDIhsn
hyIQ/fEtU/NcWMoCGWwD7j1SbDwX/y/CDyUT+C5HxMhNWp0GNuSanKrHjeygtPU1ntW3kP0FPZ6qlPyFvtQl6Z0bvupPSkv/bkE9dD0OoHKxKEvkJvgQBVryxvFtePOi
UQbwBJNpxnf/ZjqGLQrxIYHE/4HAywc8rGHEtsXVaDU3lfBU966fxE3tz0A3KweIDuC56KrGDajv8/21857rrDLSXY9ZlhaBJqbdLhUbYpzV6CUP/0vaev1LZHXNfdMH
UMC4+s9/hq6rTS6hF/R/bfvYWkHb1tsjdrZDDKD707PhFXmAbR6Le3mBWzt5QYgBAIitttPkIk5hnpag0pkYjBUrd4Rnl8wjOL9thY6XoKn1czva2+1EePY9fGQHSuY2
lltXmzjdkXVvf22BQHxrKA2nJ4HmgMhIGx4qzwg85+xozSJsv8zqvjwymne3H0zm2c8vQNNEqZgB8ohCO0Wyt50bvupPSkv/bkE9dD0OoHIl4bue74XvrBpAi/hskXB5
sOGQSaSQ+zHeSwEHDiY73UFLZyxuAKGlJHzNICuETSjKiCbRJr2HgYyrX3ljAm2I8taqJXue+34RL80Lj5h+OqHQ8Lb/521rhjLoVMECBxmtWT9XnaZs9fnizQQIPRTC
/LmdZJkur3hJ/WK+q9Wv9OYTBoE9dG5dQ9g/lyExLC90kAub32gmVtYhQArsKnOYr9QVsoJc+v+vHH8MBMv8YLkH8KjCf8rQSThdIXNlOF/FSvzN+h+6tEuvTcDDdDQh
YYMLxqQWDaCoBbBpatS7PYHE/4HAywc8rGHEtsXVaDU4t9qlNZ3UTYGFCoVwEpdKZ3dcA+iKXj4UrI7uJusdyyqUW6oMtaPasW1gUo6VMy2Ql6QO7SJoMVckaO6dVidY
2uiMLh8PrYChDc1USxmXXLPqzge+g22Bp+dJaQJvBsBTAK76n3Y9TjNbuDrsC6b6JNzQmcRV/TsBgmh8HqIb4qOXCIWBKK/SVVmNly5fYvB723H978UNd4onFOJKzv0o
kpFEAHvAxIcZJQskbG/0VtOTxHzFZjWyo5UDXqVLg0eWW1ebON2RdW9/bYFAfGsoDacngeaAyEgbHirPCDzn7GjNImy/zOq+PDKad7cfTOY+mTqIb8L5Cef35eI98+pv
O9dlglVwxFM3K97yTfzN6/29CWnvQJjzmBf7ELLbRd4aWXm63fkq42LNcTVgyZNNbymzngLMW6igjn+CMznec2bAwkPOxLg59BetQfugtp3eMVcfei6KBeqqMB+hgXW/
iHCNfMuIOZL3bUnhZ6O/J+xFzhrv4/LzHp33iNwBNE76e9G2+b6MMXPfpmcQlhwbI/bWCQyiGvDYLZpErJpEC/wK8Uv2deupdm8CKghvT/uGdKSfx23Ge5jNzT16afOt
pFOiDarTYEHmrP6vSYdqC2Ju4OJ43r/pgsYnaHd3zJJ9rZlVk9N7nA2Ol/7lLLxftmx2LvxvJJqEg8oI9mONa5W8ijBAyfcnFRsW+Pv/kjuHUTlxN25KkkkHMBxxaQFd
EOvsU6VcuOkvY2aGzayCSZwqqemhkw52qBUZoJEu63rwZiMTHZzVrZMl3f67C6wqntwWrAhNzRLdzvyuDKmnMOLD0J/OcUJ6Y8I0Y2FQ+//8CvFL9nXrqXZvAioIb0/7
O9dlglVwxFM3K97yTfzN6zH2TvHjk5joTeSqMfYw/tYTdnrdTORmuONXR+jMh6RaVZvUBWM9ISS70lT6gQOcxJszsX6G8KbWqZsktSg3k8IIeYhY/kkDOk+gnkpAP4Qp
Mw4uPdbh2w6M+fICoe0X08qIJtEmvYeBjKtfeWMCbYhqTJZpGAve3DvGd1WJKT9vTVf5cyqFajczgdCCDQvLmim8fs4B3X+3GGEtw7OQitj2Dl43NsNYFOrWQkGsrVdK
kz+nwTxmLIydUb4eBQkzh2dmgDXawhVwUEEmrgdnx33/EpVm2t5pDH+0KaXMLopdoPejuWTbTvma9Hj0YVw56R8XNw54fAT4LYcuAm4UGSOUz0sUOTld6Z949CN2nQWI
2Qvzg7IfNmS7vnC2mvFCFqYFGQRZDYjyRkpnfHHTrxuX/NWuTdrLplXpBtJwup4NuyVHdwlCtKxKaGR3htbC/ViiM/UPb8MeEeONk3N2ya9Vm9QFYz0hJLvSVPqBA5zE
26JeuBfMkN5vK7wS1VrcZQSk2CdiBWTPVsPUzbit6MzKiCbRJr2HgYyrX3ljAm2IjpPi4h/XXh+4pZBOSNhTYR5QF5vqVXi+THQ+KUL1NDLbfQNc5u9eDuZ3AtovRF10
Wxl1AC108omuYnUm2r/X74ah3rAKO5lrBGmEXif0mJbby9RFtxAhtpqCbemcyioxd5x+6dt7zHztx2SCdJFLd2Ju4OJ43r/pgsYnaHd3zJJ0QyTCX3Skojl+srRilP42
/hkmRWSlFNwJRUy/Mt0Yh4vv+0sdQ9IRSSIe0MBUl3umWd5bwkPkUa95u5qPXS3d+jSa7v5CVWfGnw6KcKE0DN+hIOssrzIM+eb8GrKMbSxFTj5AbW1ufFx8ZRuDXhUw
V6SL4/ZV4W6ltZ73M6Gq9CqeHF1/IlovLf2nzUMZH3ebdlYWl7PIqKXQ0q6FpGPpu+hz60DvV1jqZGFwsYEsiZDO506nFuxSC6t1ZhvGyGBA/UPohwg8b2pJSaPjNu12
VVoZxteUfg8lSm3Cv4KASL1Y+ejqY6P2e2GVwj5a9eeztCuflcFq9LUPtBier2SwOmZanDyVxoBgeZOAjg4DOCmO/G8ONsRIAQfXY3ibsLZVWhnG15R+DyVKbcK/goBI
vLm/xwlaTaDePr1r4kSe750bvupPSkv/bkE9dD0OoHIEEb0kFXt8aaVlSDDE1qXOy1jPIUmezd9DZe8Y5m6aSMp/biAFQnTcnlf9TCMkNzySkUQAe8DEhxklCyRsb/RW
hfvtrYwyKiJjHp3OgGe3nf41FMykoVM1f27QE703lhRW8DqghSiPwaRKdGR8cXXFN16LUwrV/ZfoBFkhaxo2D9pF5g6+kBABAL2rZHl+5rpgWdznTXbvsD+ieA5blT3q
nSSqVw8/wHqSonyLA9/sWG2oJ/a7lIGWIeClN/lfFPR8b8Od30+7/aSmg5+6oB1Dds+OSwXC1G8ofO3g7gQdlud2ddqg0chmXF0FphuutdHb9sq2WyEAh2N8vJ26EW1G
eT2/yUl6OFdMQ8D3TJxLIasmVGcg2eoWehTJ7RnsirVh9xlKj3JtCIhFC9XnqPwhlDQi4ZXw/YOriN/8ENQKWmguChAH+2iJUeWEM/XnhVypYk9vChyLjEqm6b1gNzxw
q6ya5HL7RZCRRoBuddRCCg6+rH3vdeN8Fd7Rn8fWm9eqMmpjIPJKd5qVJdjgcpX+p+5jzd59728a4fUek8rlEA8zaseLZ/Y22K8BZG8xPD3YGFklZyw8hpk6iV+Cwe46
CjNs3Ev+Y7sMVki70Jfwd7Pqzge+g22Bp+dJaQJvBsB3dhbfR4RsCERm/JbQ+MupWHnCxa4b+rffHh45yrNdgWCi/KHhdIeP7odQeocfWkWLtqx9gNQJJIePtzD3PhTy
d2dFqEswKwhzpdMZXTAk2wuKQE2NH9hwcrSgvRX2szRudrqoLwL9+/Ec01YTQUKNqyZUZyDZ6hZ6FMntGeyKtWH3GUqPcm0IiEUL1eeo/CGUNCLhlfD9g6uI3/wQ1Apa
uQKby0G85Bxr0swwc6GvyZ/mr5f0mWWxBPn8kL9Ebgbg4mwQIgybjfHbE6kS7aQTV2iyiEG4dQOp6XzlSr+6kVzzsg5NyAtJpOhm36VgeNSfm9dkCOsoACYzE494YUMK
8lfgCsN5D82qPCzHnYhi4soSJTR+IWCiof9nLXt6X5YKM2zcS/5juwxWSLvQl/B3s+rOB76DbYGn50lpAm8GwDlUFp0lrTB9DawMGCfxZxgr85cwV1ws6Lh4CevGbrVw
c77TXVikYrXHqGwVzZ0xWIvFMUFI4X+LnLyHTuriaebWimvusHDbyMQ41+dZJGia4DzWde6oFAaEJr3kj8m+1kIEm9Ya+TsJTV2yUmdvz6Lj2KSvYoMebAYY6iiN7r3P
twJavWTOLLiiGbl4vY91MBJZQpjcIYtg2ei6gWs/tQEVxXbHaM/eHh5B/25CWXlHFcV2x2jP3h4eQf9uQll5R3mQsBNt6bE9OKKN1+lvm+r/EpVm2t5pDH+0KaXMLopd
q1fM5W5WR4zfd487nSLUkYg7RRKTaK5+8RZ5+pS2G9AVxXbHaM/eHh5B/25CWXlHVuhw3M+lcTr33O+tNe9qCP8SlWba3mkMf7Qppcwuil2rV8zlblZHjN93jzudItSR
xpy8s9vSiKfmHOQR2J48yhXFdsdoz94eHkH/bkJZeUdxU0vm6hXJY7J/PL5ag9zP/xKVZtreaQx/tCmlzC6KXTcmyaTZU+RYMpqyP4dPffNlGu7cx1kBNyEXIi1G0KB/
LrDME2sRAJu5CtYzIA1wiePYpK9igx5sBhjqKI3uvc+IcTeQ9tsl6JrWI7nxfQeiEllCmNwhi2DZ6LqBaz+1ARXFdsdoz94eHkH/bkJZeUcVxXbHaM/eHh5B/25CWXlH
uzJtl7PfurrMN/BcZlQwWv8SlWba3mkMf7Qppcwuil2rV8zlblZHjN93jzudItSRoz5z82StfUkhGvFzX7JTPxXFdsdoz94eHkH/bkJZeUfz9+N1IQiYxFk+00ZOkx7J
Rnbv2attIpjNpKd49EGO6dqadBefq25zaLwuM10LiO+kYLr2ibIVh+DmScdauqDYadeVrGEPkkQ0m6+9sPfI2TA/cl1W8v7zCXmrIxO1FQzCLqX+ahBcVrRRO0Dt8Vx+
ylwBjvqCNyhzWSMXZNH+Bhanq19LzT7KjUzIrsttN1SOMFDvk8QYIBnLjEBA8+5njpPi4h/XXh+4pZBOSNhTYWzA+mGhE09VnvJZNbESy4v42oT/s0oyfFwEWPAgJ6GS
36SA37eL1ZToGcObo00xXMqIJtEmvYeBjKtfeWMCbYhqTJZpGAve3DvGd1WJKT9vF8MDYFxfG3qa0lnWkGxP6iITCr3tkdqxwulObTP5nZiGod6wCjuZawRphF4n9JiW
6+sv7N3/zEdRLHX1cYWS4uGx03VOKeCMlPVqX/daH0Cz6s4HvoNtgafnSWkCbwbAUwCu+p92PU4zW7g67Aum+rrRQfzxktIcVmiSXiwFdfbgddCXXRJpI/B/rrNz4tEI
0XqG3muFeVlsIvK5fycYsV/jMtJq6kUo3++2KGZn7ZDBuLB6OsTZMRblKTD4do8F2/bKtlshAIdjfLyduhFtRh3Qp60fFs9uOjurshYVG9q3pyAtdOyTVM4K8B83PVhF
tuNbjijgo9P8lNYy5eh/gH8Oy9zpSV7QHmQTcE6LYlL/Y2RL7Wgm4i3GewzM05ciT6YxXfu+ulC4Vy+nhkwuAIHE/4HAywc8rGHEtsXVaDUmIIqLNwgVY/+Gzu6edNJQ
UN9ebOIdEGPOlKrd2ADYarPqzge+g22Bp+dJaQJvBsD1V7kYqIesltROkhqgfSPZNRHrLUM21o9NsfQujbegpDvmDRagm2rhwFKp8j9qtv8ZPb8Cl0bUTep1SUT+p36V
QSyG2rbrcT9FYFi4DToDzDeAKq2PSdjQiYDJm00N/xNmEzfnzPYzoJL7Oj5dxgfDw+EGB1V9g7Gf+fyTH5WPlkheMM3iA+oIjFbs63LGC+u8IwmG0eIjcKlw2WuikbHa
+Z0BBHJMVShdaAOpg5UduYPDXg/oA/CBgz/cfC6gEsamwcfBesHCKP29/mTaV246GWNod+dwZN2HU9M4ZVpIYSx6Pxdkt6Vi0iSTI45OjwUG5ulJVLLe9bF7guuaciWC
JryprLDsfWvjd9IOaMsRqO+DRbQH32bW6n8EQJApXYdJeWokDOwNzREPjQnmtOICozoBmNPCbne2Zyw3KvVNTVq7JzlW2M2tfKThYkp9T9nmi+JEPg/Tl27vEMuj36iy
1opr7rBw28jEONfnWSRomqPFL+FaUfPZ+60HNcz2UwMmU2uZu3KFRZosmrwjWLtLihHFZfaNRsNdfQRbpnQULj8I1eoMWv1ywSBkTgj5Cv5acK9+Mirwp9ehgEg00JsQ
/tM6zr5L4YPfOpktF4I/bJZWP2HPEkHviDb3lJtoZPMNgziA2WtE0So55EiQTOKjp6nJO7tj6RoExqZWOiMSG9uSeKlXnelIVuLBEkWyL2JoY9EPHP3TP8Dzyshya/i6
UDfz8p1GEAopq8oVAIei6d9Gfaz49vhRSxPsZPSWZI4lQz0lLUmdXY+WlYGlNDKL2/A5nyclZyZOzr1hK1rrKVHxQVN7WuZFmQcNCEaT3iIlIgE9YV7mBazsxDh+U0/V
loczju4CjC/aNNBYXYLth11KpPN5Qdnzvigyh+N215Lo3uCEK1ydloO9cCBObVgETZ5Dd3EbNWSLbYAdddirh0lP27Y4bMAUeD0+2zJvfmfyzbTq3+8jVWk83kJER5Tt
K1nU+hFRohey+BvnzeWbHtvwOZ8nJWcmTs69YSta6ylR8UFTe1rmRZkHDQhGk94iJYF82DYLH/93rSEVsbMkdyG54+pMf3DlwQrtgy5SYH1KsSgW0x7Bb6EK5Rn/rQ8p
HmUPd1ReILbWeeDvan4sJpucyg0Ch0YAGmnQVhu4dkHPk3ZhP1y0Hl23iDuXTErLKq9PgsRSvQo4Ov8q/Z/Gze/7bYsy1HQA3kClKNzXJCIzECBZfQsrvexnx+JZEitn
A3YetUVcRYbuOkhPjxRyDARyxVWf+CtCT4SW0pdpYYPYMx4aIiz7e7ZiglK7wDz4ejiA5brjE59/dgZeNUeR4SuOpRjvSdyXAuB3T4M7ZyHVY5LSjRTE0VUwi0575SOo
aIAT+6h2/ykPNL9POFEc6tMGDAUmC3w7QePi1qNifadNnkN3cRs1ZIttgB112KuHOphwATLtaA5C0EoIoK1V9IDkJJ3LKg3L5jDZrCliWAknycArXlCYlBQeiHAsCVvw
JDqMbhyQNYUeGZPGvOtNKXEsTeAHw3T6CXj5P3XgVhdN31NwfuplLS5k18eIh3MZd0+xhQYcsTXEWBilAkM+OqjN1RLs1/jxqLyQWUJDHXoccvEASIrK6a1Gb7vYbGKJ
m5zKDQKHRgAaadBWG7h2QTg0Ad8bHTH0O9V5v3Ii0s3o3uCEK1ydloO9cCBObVgETZ5Dd3EbNWSLbYAdddirhzqYcAEy7WgOQtBKCKCtVfT4VaHtx0CkYlxQP6Xl1eAP
aGPRDxz90z/A88rIcmv4uvLBwaWK6KzhUrndNm2ahmffOzaawqgiGoUD1xd2TGF/coviJ1STxZvtHQsINp7UrG/WUoMdI8CDkzmFhti+E25svRpsQjditODHq882n+yw
bg4H6JiYSC/O80axpbXvYwN2HrVFXEWG7jpIT48UcgxFUKVbvvvLZZ/KJMccU0X4uLXLZFiCUDaKOO4X1VM8khvcy1L2oh52NuN1jEIGP9PDThk0HSbbuy/SuJkQkbxp
htPW1liygKfyLRlWMPNqvWhj0Q8c/dM/wPPKyHJr+LrywcGliuis4VK53TZtmoZnXqKbnBlbDTQNTHhHrFX/7DGKar66mO5F92y6M4r3c2XS15y4dWbUQPIt4bNC2dHB
Ck1+Y6Vxga5grwEePdkXDyI8iiJXm0omLsIoOrWYZu1R8UFTe1rmRZkHDQhGk94ilXjilKBCU7nfLdO2gOCvIfTybedozIXlttWvTsVAQbMnQTz9xdcXxUAGpPSl5tXF
gbC+sAvVyoj76rFVThQEJ9CRtu5cMCfNKZZ9SFKlc+n+ANivyuroC0T3qa1vste3Gob5YmFL7hv1iFQGg7XMzAlrWl5pakOuXirdKUI0qGzNbJWwNWUNCLEsoiOSlAwX
+JBpn4/idodXrgcaIILfuHRXEZHINZU8XBllCnQLdjPokUkWG3XA7NJXyPFvx2JjMWKOx8A5xOmmWGCUVl6ZUZma0cBnaRqHeATiaOiMOfAjJeAVDaZNQo0ZKDexHJHL
u5xlB1pxWIR6CuppDaTs5LDhkEmkkPsx3ksBBw4mO91BS2csbgChpSR8zSArhE0oVNKB9ZHwR+ci0XGrbYSFHwcimKGPvF8h7U9eA/KR4boxRfFLDC2l0K591q03nmxD
BwIX+vefl/HuEIrThqnl35IqXtnemfAt+JjJ0HF/SyKVTMKcF5CyZ28wV8cknzvF5yFuAjkA7rlyLgNpfI8TqS36RSEeHNUdS7mVvlbeHova0fy5lDxJelrN2dsTeN9N
HjioZB9pk/x/C9OSAXDRAqYb16riLI8lJCSLuLATS1e/8VQFzGdOqu9R6gRvPJo76Isoaq16o+JZhpMyTRtQulygoDDDXIPrckRsCfvz3tQnmbo0SN6wfiAkjK2z8qgn
BTJ4anjRwm9/QMN+Vb8As6ME8KihGeeHTCBcge+3AtdQHssXyJcGurlboe6713mH1prcuRz/tS10bllV+/Yaz1G8ALJjXz2FQZ93P8eMAo6CBg4dyqGsD4BrLCozQI71
+z9uuJYMGqrqaF32wedOqd0q9JGdi89VfxM6JuX46xz2Ho7Rsb2GAAFJHQ/lkqjFq19ONxYjI6Zijxu244TMdgOJX2gtMdr4/ZB6xXU/iHkBxO8XyDCigwqYoCu/mbTw
d9dBHMqvmHh2/EmWtxS3NKfA37fEVK7/SLks9VNL7iQxYo7HwDnE6aZYYJRWXplRdfAGlYkYyVDo74KFq6wkSmFz3CvuUG1cAHCKe8eTWABU0oH1kfBH5yLRcatthIUf
OqH9u0jx+x3skqzjvcgwa8wvMa7ShBBvGMt9c9aKqRCtS8Rk0n0EhJ0wTqO7J9CoCZmyJj/YMtMCuiYhR2YvcRIkWC+iYfxPA2Ci+ML6Mr3LDbdYjm5I2xmIzE57bFRE
pj0UI0esNg5z/ZE4wJ/jL/pJw6C1B3HcpFI+6zVjYydRhF2qD021tJd/pRKmvYMKSJ4u5+7zNgEscFF0wRfpMviQaZ+P4naHV64HGiCC37i+I4+1qTaLVFRmspr2/8wg
dmjknOfpyrJ0pNw7TPc4sPQo+UZTUKGwTHAuiBE9LufVVYHaBVoMf32Ufwty0BzC84xt+d57sD3dAxzSuZEu3I1sZWZafNqzqrqnGgBVQFJHDgYTvM6pZ8uDwmH/lUhy
WQNREHA33fYbU4zfhci1RsuMcA8R83ylGp4CdWFdv/O+pnNTkmhtnr7zRuckaS0Gukg35KcnVn2Sxv6xt5aCBL/jX/CAO7Zaik6mU8EaU48dUXoDeJAV9q3aWAK9bz9K
ncsMjweEuTQFpG5np54wUL865IZRJ99YfRr/f3NQ7sdZGrcpv7/N6uDd5rF4Rb2Fs+lLC2hgQ66UK99IMQy0C5dcGboysyaej6VfpR+DxaxvzbeLIaTOYWowhlUNoagg
/dBjI+Ab+dO9T8e8q80Vee3qZZISEP5ZcLbrkcyEmgW0fw09k64WYrOi3UhCMo0tADfedmqSGqsc7LroeGb7hYws9T41aO9l5MDGSoIRtRDAyriLsjDnkM+LnQAKE6/e
zmMOA+e1hTpmDMWl8xWKsWps5F3r4/eOJ5IYPdA+DH/+qMh1nuK8FjazyxiFTwI2y+wU5QXN0cCIv+MWOYck0QJgo8PZzCXV4UWMiFKH2rJNPa2n15V0mmGsetuCf0bI
54V1JFD3FxL10jWzAMCR37/935kGSVvgjxEIcZc9QPOEJ6pM2Q6Ljfp3WvXo55yewWBMIAjyiRwFSbQnnzNuTLBMGfIuzqa4w7/taFP1jMxLh/v7/t11t3koRf+jMbbM
Ilqz8oBZkfxPh2clIKQXdbEjJ7dxV56wv0cnrw5qdtTpzKbZ1a6H4+3stoxE1k5Whubch2BapsRhVJFV6YMH6n4vL0x+qaq6jNrpf+G+gQkBuMFHGXOV/+W+hgYvjvau
vsW5kfrNCNenQLpYAwyePKfxkbO680bd5yKQGoxvVVBg5KxpumxBpTZVX5UYFx851SmXW52x0rxAa6u6iIeYu4+TSZa2RuLVbgc6irYm/cw5LCEdyCFLULoD/2ZNzwLX
ixP/i8KkjrgqT1x/ZxWD8wuFK2kox2n6XEJRwjMpBc7j/VWDrjgEJRUfGZtQsAoruCrdV4WsUfq7MwgLe3d/uNCo5MKlboVlRIWPCsagzADuCj0kJOWIodP4rbfaj1p4
BLGnT6SSIj623sX3j6CWmEPyWKH1CKIWfsqpaEGnl89TtZubFmUBuOtrtmpc/9oaaAvqb6yu1N7OQYhs2sq91dYJ5UPb5CrDQRbD+Vt6RTxrJDURTMeQFoXZ/TeccdxM
AdIEtGFZFuaDNyP6a+2bOZm4WkY6nwoMrpor5Mrn2q/dN0uQrQ0RdRHOwEuOPLqQddNeX/Afw8Bi4succlByGMwl3bru22/lIOFZxLRLTp6fgFMR3Qm+9cJce9y2hGAo
Xyf4B+Ggo6Bg9ZDb9dt8yYCqKOqhxwprYFUFnjz5pQl0LC9ODWtHUAY9oSg8zCXs7go9JCTliKHT+K232o9aeGm2J6Kqosni0JgodfpGejTDwjqHCbs5p+/aMc5XMh/6
GQ6FZQ9W6nleUpbDzuwqZTgFs9TUgk1J8gnsVRMp4YiGod6wCjuZawRphF4n9JiWVLtOBSFPTuSVSuWE53RV4nIC8UjYT96taOuFkw92gJDEP/alIUMPgEscyvycoPkH
Y8M7UCss/vJoEobUATZzDL7FuZH6zQjXp0C6WAMMnjwjQHRnoZEX6XeCkn+tLYoycVpyGETzDbpavnrwiM7qO/FhqXAGdR2ppjNTAfXnjXOjE0fUSkXfAOyoRQHc0uVl
jJ7UhJ1XSEpxHrlf6J+4yPcFXzd1pAKGsnsT8XdAKonj/VWDrjgEJRUfGZtQsAorMA8l55K/ot5KUmSk9hBsmxMdcYXoZrdJlyD4wYef0lrHvWdXoiVCTUjBDLYW+smq
6FwXxquMBv0Qb/QOZzOaMqaGlhsErD1ydQUh1bs5a8Jm96E8/OO/ECafThQnVV/8z9K52jyr9PY9MY+ZxL+CjlSpZAjU7ti0xL+BuF/KCcj5ayVTXu4H/7gJtehdCOJ2
A8v4x75/toSmOAVI0QnOxZv6mg881g3p/GAsr9prbWOGod6wCjuZawRphF4n9JiWVLtOBSFPTuSVSuWE53RV4nIC8UjYT96taOuFkw92gJBYC5P2KXXdXn4D98/B49Hi
11gTaLpje2/e16TRhUenY+sWpPWXAKzPguLaP392iAY7dZOF8i+SFH56YP1tVJL0poeGgE3TWSqHzRSaUkGSkR/ZLzIbE/o5tIwYrSn3k0VM+C7TvQzy3uLaZbmN3QgW
Sa2S6Lwz0LdVPOHT3ud9NQjp1539lrmXWa4kgn74lVsS8IDjaqTIjwPY5bN2dWdRYUxyYCtPL/PCedC5ivOUfUjfkYrw9r2IJPA+SLFkT2x3/KMBu/hlBGW4vDv5UnEa
1XsdR/L4QB3uA8oRNw1RGIwmiAII/9vjEj+O8rHqIMEiKI4grLzGmCC3apA9NuUggcT/gcDLBzysYcS2xdVoNY+VrqYJafgeSwXlloVXgVySbEanb1EvQZzEMMGLD0r1
fw7L3OlJXtAeZBNwTotiUmRfDGzIEUoGmkY5KymTiQl0ticFDfZCAbR3cp5TKoj4eraMep6T5+iQeNZY9KMyu00EUPHXg8757JO2Ok8C73DhFXmAbR6Le3mBWzt5QYgB
pOTJ2Y58cA5L+4e0Y+9Bl95xAcN/8yzkabJ85efgOeoW4m/y8OwvBW1NvM874JKImAPwB1O6PioAuCpB7ynDQH8JoLRnZqMe6vBK0qhm+WVB8BGr7Rkl53LMxbkF8mbd
BUsdlkP5SAKfpZMCzoYQyAzuIM06pzpbRXiJLv26XKexXKrry+cnusk5Ft1Rx3cxSNp/bq2RGTNMZ4VMATmv7aKN9h7/YrhMNzy+x2UbrIi7JUd3CUK0rEpoZHeG1sL9
WKIz9Q9vwx4R442Tc3bJr38Oy9zpSV7QHmQTcE6LYlKl9EEVZygYBSOV8ZV44oJPlQHQ0yeg6C+2+8nqTdQfjNVR60TO3viFWeKmZJbotYyWW1ebON2RdW9/bYFAfGso
mtCxprfhn08DVStAHiC/IPoFcK8jx+fvKXUCdGNQuDjDYnATX5hm9SJeQskwpJfgQdXIX3Sn1wmtxel8j6zJuaQlsnjusIuBIgyZcdiTt/7/3EntTVht+LFYJyMfS/In
c+7upI7xFTlX7jsDx4Qr8UN2+mdVY43DgeGvHCviGAHvxYb6v85XaNRq1clLeo33AraCG6rOiVuo0XAAE3BMHn8Oy9zpSV7QHmQTcE6LYlKqx/a91VAIfuLhzgveArwu
roWLutZrKAUX2ZbmpZJspA8Ebg8sz13Q8DQwmH9cBYsGHgA2uxj8T+QNpUDmUGaGyogm0Sa9h4GMq195YwJtiGKrTJrjigGZf8ZOg6zpjRliq0ya44oBmX/GToOs6Y0Z
bSHsar1Srnt8N+LjBvGRkfG9Kqkoxg4HFe+4g8ZlLHTLr2uNg5FcPXwGqSyyL79tTCDFG7YozWp/1i4mXyP+FhvEmR5+qYjjS7XnIhwpagripH04BJdhWGpGeLx3Z9bh
zGtqE9C9UB+KCTv0Dg3Gj9u/NzR+aSpJ78VyePbcEVOh9ksNzna/Hu0lkyltEJq+WYT5ugrCfswhy2jRXS9aG18L3p3I7KKFLCjMOSsozO9GKaTpzCHzuuTDMbzAOGwm
FSB6SQ+dtAc6Yntp4OD1qV4PhBM0ItUSvkvcEL9cj7yGBvf7F0OZDvXHp8Zvki1F1ziIKB76JJCLvrs9HVe4De6/zB0MxYOxK1Eny4B67OanjHXr8ONHafV2lAQeRpdL
tgh/zGnT9lwiQk4qBGWWAoR0kbPeQHVTgE8feqlLdLq8n3igUvTgJq9rvcScR00O7c7a7lt5P1BcEpYf+MWleE+uTFdqbWfPE3VgKOG+5lvEJwB6KgmeNGdmM60Yx6eo
K1/jf6cxlFFSvuEDkz5mbUwgxRu2KM1qf9YuJl8j/hYbxJkefqmI40u15yIcKWoK4qR9OASXYVhqRni8d2fW4cxrahPQvVAfigk79A4Nxo9Dl2PUnmVD6WlF8WqNq5oi
PI4reyvlw9cnLb95OxAhsR2DmxazdVYRrm8aekUXrVxptieiqqLJ4tCYKHX6Rno0++p7LVCnzp2bUNSjZhzNUwJW2AJKxkzQkJBOGlfO3/Zqs8qIPIuRYfmUxuVREOXr
shJlfCLdQMmV9nJR85F/RL99a47u2Raxd/DB/5JFI6Q8AHb+Q2VZHXZxQwFOY9TW9iB338VMTSltF4jjK7J4ljdg+x4zYpJBkVyAN8IYCocFY6L0fAe7rfVxffpEASr4
x2P7LejYNCkCfcbc/pDjWcqpOD4iocFQfULBOLcR08AyJX8ezLtHBUkPcW28LjF+H5UVdLHDE9vrOK3XfFZNwOm2Q+/OpZ2P7NCqzfp9om0f1ICbmf5o1/vqVfenaUk2
e2+ZRdxYl6JUY9tCTd8l2PaeYMyWR19nt/1HEY5EHNp0v3xlgo96rrRfsnvFczm/4PRdbGd4125LX1vPnwYNe9PsoPW6wGQ5WBqkfmDE0QyIL2Qrllzq7oZ1+3/zGlcx
r4e+6DhhkYnv9zNSxPjDkJezNjj0XmKI7f/5+BLp6lr/jGcs50RVbo3kY0IjN8hlli/FN1TnLwVSCmr2UehsmWIPVAn5h4SAfxqlG0tevWhrrB9Ab9opTWmFVy9ySOwM
ifU8OATdrY9wNC9P26f8K2vceNwHkOhnb2aNaAsaA91hKRmh/hBb114zswOPouJ2nN6N2+Zj1U0SdMaEfxlRKgz/802+kTEtjYgS9J87MUEl/WCBaltqbOxgnecFy0HR
xxl2PqibvuTjT8OaGjn3iuVRmVJM2MT0jSpTRy52J/pUCs4XIPpWE5LmkkUGtGtNy1jPIUmezd9DZe8Y5m6aSPE1bJUjCHo8ds3hjCZLFpjyBwCwFKqqhMxUO80gmGxS
GTRWlTJHuSNtvjqjD0OVnxdVbJ+AInYJYdwWo8+KBODHyxLlHY9l9cWJNWOK+NmcV2jv7ZmVX1F8oTE2wFuBPaT69feX57FABo8EaWxYNY/FSvzN+h+6tEuvTcDDdDQh
YYMLxqQWDaCoBbBpatS7PVosW3UCXQQk3RlLOknwdd0p4Y1rwkGql8hhdDbM3UG9x1/doDpqWQbO1tBSDjRwXVPmHDo4vsJBaslb9LpaHDhA5phuOwivLCMzJdXbfrY6
j95ZbKk4SBaXBUh/KbbzTfSmD+v/l6r3tm+FeyQirncbFe6HWHX+cTyLBFBP+I/D0d1psf/xfWc/TWpQ7tZJE8KUVd6FplxFJsJO/5iEdn+jDouIZUCh3l7Nw71+vSWz
TCDFG7YozWp/1i4mXyP+Ft3yYHWWN8D6p6lcWJN6YlCXszY49F5iiO3/+fgS6epaNbOvmCrqAVCLJhg2nOyIqnRuTW9wDk/IReMqU/gcG/lsW6vHpLfb0FxF4Lyh9Etd
xpVdUBXUwY0NyJEcQ+4LTVPmHDo4vsJBaslb9LpaHDgf1ICbmf5o1/vqVfenaUk2e2+ZRdxYl6JUY9tCTd8l2PaeYMyWR19nt/1HEY5EHNp0v3xlgo96rrRfsnvFczm/
7sekIUeySsZ2vQNfhjLEs9w/Dxs7QlTAd3WebNRkcjNe3A8pSai6BjBtWRs69CTg7B3gNiwmYPIM2+/wrPPjA5zejdvmY9VNEnTGhH8ZUSrmTBrc7KXnZ9qY5KBOM3xs
2I6IELSJzooYPVc0uysreBHRCf+sWOv/VlpWLLcN6Ugw6/WrnVkocg3MOirOcjv7/AHXG+3jONGvMOd0D7ysl2K5p3oljeEF9Pi/Iw6/qY55Pb/JSXo4V0xDwPdMnEsh
ovmqbUBmgA3ycVX5Kqb62DG2uoc16NEo0HgOljidBS2gKL9NkOckOAnPlY2Yjh8+iH4WLV5F57C2+TqA7g8UZHMx99rPIMRQpxP8oki3WxLvIYP/ClSaUuTkSbnUlQAH
RUVp4dcA/Y0fdoDZ5Dp69kZHncROMzshjNQtH3XdrNUzTPz38Hte4HN2x5Uma8TKqjJqYyDySnealSXY4HKV/oUvc9veQDEAR6qgKRI5AOgJNyZIv07XoXPFpwTctzei
zFbzN6wAsXdChYNnYMJmadmY8J993AVo0sALQqAW4NK0ad01QHD/L/wkU17k9GNIAIitttPkIk5hnpag0pkYjBUrd4Rnl8wjOL9thY6XoKn1czva2+1EePY9fGQHSuY2
0zxcTo8fEbtcGyjeqzEBM5FYdNXHKaUrTznGZkq88h8lENJC9xsUeyGkMai+uhRz2dxrq7jm2HM9mNpIUqu8ikTOuYLZarIiS2jnSeYtIwcR7LVfB+cIGrCxYMULpemx
6+qfd3CPWQcEPXt5+WUf4jNM/Pfwe17gc3bHlSZrxMqqMmpjIPJKd5qVJdjgcpX+l/FHLkqUmNBGZmgSe+vjACGBqMp/cNoIwlE6lUGtdWKb1d30fhZdEfHJbM4Oho2H
D+W173FA44+ij9jLt03Cu5uIHW7Woqy8NwsMsOLIjPBZhPm6CsJ+zCHLaNFdL1obXwvencjsooUsKMw5KyjM70YppOnMIfO65MMxvMA4bCYVIHpJD520Bzpie2ng4PWp
FQ96AzJTvBQyuqy+dlSWz6m7sKC3KzBBmrttERJkCa7aQbnynrv7LxzVpyfafmd2e7WisVj/ml81p8mxu5NXBUvUYVGSemEABXG3Alo8710AiK220+QiTmGelqDSmRiM
FSt3hGeXzCM4v22FjpegqfVzO9rb7UR49j18ZAdK5jbTPFxOjx8Ru1wbKN6rMQEziQPyUnORoSSgGE5fkqMD2lINTer3Kz0TWXVG+o8BDEoLKJ+irPbPdcovKncP6oO+
1gZq+5jr9rlsALHTGfToEMVK/M36H7q0S69NwMN0NCFhgwvGpBYNoKgFsGlq1Ls9OpvoGAam1gfhSKUiz/ebrZ6S8f22MAmXsYnEn3qTrk3f/vdWrYWl8mQuoqlb3TJN
XdmI8kTqGVzr3HrN+/3Rsah58vqF9js3jYDkPIZLDBdlGu7cx1kBNyEXIi1G0KB/LrDME2sRAJu5CtYzIA1wib1dkS5SE9HTHnz61lKxvFFES/notpvPCg7EGoG5ASuj
jML2jQH/CpclN0vzx2jxqgson6Ks9s91yi8qdw/qg76h5penjg3uzTwziKM9XB0wZRru3MdZATchFyItRtCgfy6wzBNrEQCbuQrWMyANcIlI3eaN0pwarTNl7XbhhYEH
/vym1PBV2F4nOYdsXBY+YTrCnGWJYzXQ57yccw9YPH6lyUn3r3hkWqQPp2ifG7toRUVp4dcA/Y0fdoDZ5Dp69qusmuRy+0WQkUaAbnXUQgoCVtgCSsZM0JCQThpXzt/2
0I5inK0eDCBMfS1LYITJQoz++dRTErPjK3GLYFlEFJN8trMPEc3qyjdk7HjIO9Zvw20ADCmedAEM8YbEjm8siKOYwGG34kuoZmZG8S5uVEFiuad6JY3hBfT4vyMOv6mO
55QaPRKxKXzCC+ylBDHl5M9uymSsJPCShBysQLR+tdKJ+bjlXRNr5Mu4Kt8mlagCEVhlipAteiQVvGTVOFkw624JjOjVfPcnl5tZi14UzgRhp4R8xKBpxk216KVHUoq5
H9SAm5n+aNf76lX3p2lJNntvmUXcWJeiVGPbQk3fJdj2nmDMlkdfZ7f9RxGORBzadL98ZYKPeq60X7J7xXM5v5md1Af1ktoQkvymFo0DKbwnzTqbIdOOhw1Qy0K44qo5
YrmneiWN4QX0+L8jDr+pjnk9v8lJejhXTEPA90ycSyGi+aptQGaADfJxVfkqpvrYMba6hzXo0SjQeA6WOJ0FLYJAmiy8Tx2m/yyDOP9doZ4GP6JSTRAS8yD4smFcCDAh
iC9kK5Zc6u6Gdft/8xpXMevqn3dwj1kHBD17efllH+IzTPz38Hte4HN2x5Uma8TKqjJqYyDySnealSXY4HKV/pfxRy5KlJjQRmZoEnvr4wCpH81Ya0YNEgWG6x/BGgor
rVXWP4rtvn/TeB4C/VcbtMkPxshis6k3wBai0mSn7IsoUcO/GVp2UFXJ+3r8zHni9p5gzJZHX2e3/UcRjkQc2hvCv6rUSrH863tWp5+0xN7SJY7rpQT3nIHj+Ix/+aR7
f6XnZ+BrMBMZySbSunqlVCoaLAFkERvzY7BR8z4oKPWoefL6hfY7N42A5DyGSwwXZRru3MdZATchFyItRtCgfy6wzBNrEQCbuQrWMyANcIm9XZEuUhPR0x58+tZSsbxR
aS4fxcEZGpZJz5wYw0Us+0gmA+h8yut6IwK1GDJEl99iuad6JY3hBfT4vyMOv6mO55QaPRKxKXzCC+ylBDHl5M9uymSsJPCShBysQLR+tdKJ+bjlXRNr5Mu4Kt8mlagC
ESlrRNN4tFx6po4ixf+RZolpfx+izkHqemI/e0eE/D4/nRiMkyRLSc+NfEaC0O3U8nL9WLxkqIcqYysWNB0WOAVjovR8B7ut9XF9+kQBKvjHY/st6Ng0KQJ9xtz+kONZ
Ye9YKwduGZrQiyfzHq8vUc/OikCYPLoJ4j+sYgB1JN2AINnp5+2OQP2J9ch25ruYYrmneiWN4QX0+L8jDr+pjueUGj0SsSl8wgvspQQx5eTPbspkrCTwkoQcrEC0frXS
ifm45V0Ta+TLuCrfJpWoAhEpa0TTeLRceqaOIsX/kWZJ83ZILI+NlQDPaMObJaTRXw+0u568u9A15ziOPOlliNTZ1OBRvQJRRKkI5NZHT1ih5penjg3uzTwziKM9XB0w
ZRru3MdZATchFyItRtCgfy6wzBNrEQCbuQrWMyANcIlI3eaN0pwarTNl7XbhhYEHLd50cE3gDCD9DMmHwcIt0eAmkVWyvcvkoXGufAE4sB0wFl4NW9heg8WvJrfV6jcK
cXUrvlAL0VoCjylYnBvXhVbwOqCFKI/BpEp0ZHxxdcVBS2csbgChpSR8zSArhE0oUZVEAxlAQp09j13XdbO+0Wpii4HdjP6f9fW8zN9yjy2uv8699+aAStIUOd30W+PN
TCDFG7YozWp/1i4mXyP+FhvEmR5+qYjjS7XnIhwpagripH04BJdhWGpGeLx3Z9bhzGtqE9C9UB+KCTv0Dg3Gj0OXY9SeZUPpaUXxao2rmiLTt82HULHyNyPOgm9mfKF4
TfpleAfwRZ48V10ufVjzrFQKzhcg+lYTkuaSRQa0a03LWM8hSZ7N30Nl7xjmbppI8TVslSMIejx2zeGMJksWmPIHALAUqqqEzFQ7zSCYbFKHUenT5V3URibkcSIx/gIJ
g7EInUnSRJhweTgfEE0YnUDmmG47CK8sIzMl1dt+tjqP3llsqThIFpcFSH8ptvNN9KYP6/+Xqve2b4V7JCKudxsV7odYdf5xPIsEUE/4j8MGhynygVufI9lYU0xur/vi
ec0JLmDT9NfWyTiMfb8r+2vceNwHkOhnb2aNaAsaA91hKRmh/hBb114zswOPouJ2nN6N2+Zj1U0SdMaEfxlRKgz/802+kTEtjYgS9J87MUHN8E2dM4Y/mo4JmHWwVplU
PIfD1a93Dx9SxC0X+BdWVEVFaeHXAP2NH3aA2eQ6evarrJrkcvtFkJFGgG511EIKAlbYAkrGTNCQkE4aV87f9tCOYpytHgwgTH0tS2CEyUKM/vnUUxKz4ytxi2BZRBST
vMeNNU92mUUtObYrLMkCnWK5p3oljeEF9Pi/Iw6/qY7nlBo9ErEpfMIL7KUEMeXkz27KZKwk8JKEHKxAtH610on5uOVdE2vky7gq3yaVqAIV5GJd23b5YfJJknlcEaP7
4+QMCyIDwNMC6yu1hC1JO17cDylJqLoGMG1ZGzr0JODsHeA2LCZg8gzb7/Cs8+MDnN6N2+Zj1U0SdMaEfxlRKuZMGtzspedn2pjkoE4zfGzwPVzNTzgqIiLUdVXETVX6
mh2Qj4YvZnGvpo456oWECDZvtuZJYR0gyILRYvpEcEc5853KbggZp643OPjjER6rAIitttPkIk5hnpag0pkYjBUrd4Rnl8wjOL9thY6XoKn1czva2+1EePY9fGQHSuY2
0zxcTo8fEbtcGyjeqzEBMy5TB33nGvZNdmWCRSeKEcAQJz/PORypRBSAM1lwFXCJcXUrvlAL0VoCjylYnBvXhVbwOqCFKI/BpEp0ZHxxdcVBS2csbgChpSR8zSArhE0o
UZVEAxlAQp09j13XdbO+0Rgqv7gW4u8SEFchZHIJBeMbE2Fy09tu3YCupcBSfUDTYrmneiWN4QX0+L8jDr+pjueUGj0SsSl8wgvspQQx5eTPbspkrCTwkoQcrEC0frXS
ifm45V0Ta+TLuCrfJpWoAmn34a9o+aBqO9ZOjoBc96hM00/RSN9RhfomrF8iwc4qCRwALsl83lawBCLfERBtZBo14cbmP9Os+H2Q0v/TytTGwASgfC16ZKW84zpDmgE0
cXUrvlAL0VoCjylYnBvXhVbwOqCFKI/BpEp0ZHxxdcVBS2csbgChpSR8zSArhE0oUZVEAxlAQp09j13XdbO+0X0V+Irb4F8E1sNaTgxqWRjvKIaFexgGbjgzFPkNDvQd
8ISuyG/xNGUsL68HC8PVS/uRQhLDr/SwzknqvNs6CygAiK220+QiTmGelqDSmRiMFSt3hGeXzCM4v22FjpegqfVzO9rb7UR49j18ZAdK5jbTPFxOjx8Ru1wbKN6rMQEz
I6RxHNwmt62zt4XXA0KVCibv8m362gBvnRlXyoJzUK4Ag+KYT8r8hfVAKNs0HKaWRUVp4dcA/Y0fdoDZ5Dp69qusmuRy+0WQkUaAbnXUQgoCVtgCSsZM0JCQThpXzt/2
0I5inK0eDCBMfS1LYITJQoz++dRTErPjK3GLYFlEFJNpW1Wgs9nt8xsp8HhXjp7818hNGCBSwKpQk2D5HTqRB2K5p3oljeEF9Pi/Iw6/qY55Pb/JSXo4V0xDwPdMnEsh
ovmqbUBmgA3ycVX5Kqb62DG2uoc16NEo0HgOljidBS20ypEzaBRfPkIu23JUQHiYJK04MaXLnpP7xdDGSwTNHScKqk/vbN+BYEfr71rodWoOlXWy0OmPXpKH+eVrmqiH
YrmneiWN4QX0+L8jDr+pjqK2thRXLThPFCt8I6GwjekCVtgCSsZM0JCQThpXzt/2e6uYEDGBCeB6jVOmJepGO8xgyYbQfwpsr7CPZ+zTwEkd8CJcJNbOv3xagkZAXITi
6IBT3spaPTZHNLpLoH0b3vBJd+ZYYhAvQCWoMynYfwulEKSPnnIOOwjcjxZaAwbKr4e+6DhhkYnv9zNSxPjDkJezNjj0XmKI7f/5+BLp6lr/jGcs50RVbo3kY0IjN8hl
li/FN1TnLwVSCmr2UehsmX/BIcq/yYOuS+HmorWfN1AHtb69EprGi7Q2/yHK/chEYrmneiWN4QX0+L8jDr+pjqK2thRXLThPFCt8I6GwjekCVtgCSsZM0JCQThpXzt/2
e6uYEDGBCeB6jVOmJepGO8xgyYbQfwpsr7CPZ+zTwEmNlvMc5O9kDDU+Y1rOtHHaI3kIkn+V+cb+BUi80/Y/f0wgxRu2KM1qf9YuJl8j/hbg4mwQIgybjfHbE6kS7aQT
z27KZKwk8JKEHKxAtH610qOrrqDordkDEZB/8XS8tdh9hRCDvhg8T95i00/2AvQbmyur/+25BuZHWskRmqAGrFfYqMQyXSpaYaTTDf8AVbBptieiqqLJ4tCYKHX6Rno0
++p7LVCnzp2bUNSjZhzNUwJW2AJKxkzQkJBOGlfO3/Zqs8qIPIuRYfmUxuVREOXrshJlfCLdQMmV9nJR85F/RGB0tdb7NAk4CmiKwstw8H7R9aceeJe1GcQGQ8dLgzEA
QOaYbjsIrywjMyXV2362Oo/eWWypOEgWlwVIfym28030pg/r/5eq97ZvhXskIq53GxXuh1h1/nE8iwRQT/iPw7Vwajriimhd9Fd6e8ii79vzo/3Kt/paUxNAH7Dfv5Sn
abYnoqqiyeLQmCh1+kZ6NPvqey1Qp86dm1DUo2YczVMCVtgCSsZM0JCQThpXzt/2arPKiDyLkWH5lMblURDl67ISZXwi3UDJlfZyUfORf0QsVnnrxBRfsHb/VklVrA9j
NFO4Pd6Pe9/iQrcCw+nUeUDmmG47CK8sIzMl1dt+tjqP3llsqThIFpcFSH8ptvNN9KYP6/+Xqve2b4V7JCKudxsV7odYdf5xPIsEUE/4j8PxCQd1GPx5pBZWUISd6cd/
CxSXL8NxzVrJGbaYA/PJ+Wm2J6Kqosni0JgodfpGejS5B/Cown/K0Ek4XSFzZThfxUr8zfofurRLr03Aw3Q0IWGDC8akFg2gqAWwaWrUuz2N/X9LXEoYSC6wgLxklHRl
dwqe4SWFm1Il+yWCYkd+Nlet4pL8OkwkssjWE8wXwuQxMQse+3gBOHJK+stqzc5UuQKby0G85Bxr0swwc6GvyZzejdvmY9VNEnTGhH8ZUSraroP1ewkmSE5B7ceCkiB4
QVdrrygfa/JsjE8BDMrPh1E3FCA53B/6xh0J6oLQi6Xz7XZu6zv0u6wl5BnlT06au5xlB1pxWIR6CuppDaTs5LDhkEmkkPsx3ksBBw4mO91BS2csbgChpSR8zSArhE0o
tuVCcGW32kAlAuhO13mxO2NqLmcmjwUzidisZRCLF3izXIDX04vNFlezOT3R+KtTpbYcb7n58mz4Zl2so0+dFjExCx77eAE4ckr6y2rNzlTuv8wdDMWDsStRJ8uAeuzm
4qR9OASXYVhqRni8d2fW4Sn/FIfUPfdjBcn/wS4a94dvf+NaBIJkC4UO8SJcWxdjUgHrG25+iNLGIYcycrvwnImfrjMnlhYLwXmtj1/Wm2rRNkbEmdQiZ8syHtUMyblk
Hz4JQB3AqneLRRmUoeflBUYppOnMIfO65MMxvMA4bCYVIHpJD520Bzpie2ng4PWpIU9vQaT01+J/6uaM/ESMF8secVvkCCK9AocRHnHI7JhRMkyWM9YkJ4Xn9YFMLg/q
uatOmFl8qxWNkimlnOK/T0VFaeHXAP2NH3aA2eQ6evarrJrkcvtFkJFGgG511EIKAlbYAkrGTNCQkE4aV87f9mqzyog8i5Fh+ZTG5VEQ5etp15WsYQ+SRDSbr72w98jZ
Q/jL76RbHK8IKr4WGYg4+jGz/+Ggnzm/qF7Q5dI/3QHLxwsG4enYdRl6rcF76nGx16zMKTOz0KyjZjLdTDLU7KHml6eODe7NPDOIoz1cHTBlGu7cx1kBNyEXIi1G0KB/
LrDME2sRAJu5CtYzIA1wiTeGyw+b9QU9jBX4TgIhauj2lsilykaIDA4W1CkPtOPP6tntAx+uiwclYt8n9UFrZ8KgYk5xGncPCk/kBlA6ew+VGnuFL3Mq1GP9nf5unVIG
cwa2z694vnjnR6J5cGSkfFVaGcbXlH4PJUptwr+CgEj0pg/r/5eq97ZvhXskIq5336Eg6yyvMgz55vwasoxtLJSd4xqF5zB224+/OnAgMEpQdhP3bENU19obsR/j4KiK
NuPiF73enmL3njksge7sn4dbC5eUnd7oBOiM0hzniIxe3A8pSai6BjBtWRs69CTg7B3gNiwmYPIM2+/wrPPjA5zejdvmY9VNEnTGhH8ZUSraroP1ewkmSE5B7ceCkiB4
6/xv1liDGd6SPoy2YIMt9/A2jtv9rMhTWtdlYA6C4WxRMkyWM9YkJ4Xn9YFMLg/qtfgJPaNmw4kaXaD5PgbcDEVFaeHXAP2NH3aA2eQ6evarrJrkcvtFkJFGgG511EIK
AlbYAkrGTNCQkE4aV87f9mqzyog8i5Fh+ZTG5VEQ5etp15WsYQ+SRDSbr72w98jZG3BbxZDYFjr/6vzxFFoW+zGz/+Ggnzm/qF7Q5dI/3QHLxwsG4enYdRl6rcF76nGx
hcVG00FgUgzIOn/rD65CUKHml6eODe7NPDOIoz1cHTBlGu7cx1kBNyEXIi1G0KB/LrDME2sRAJu5CtYzIA1wiTeGyw+b9QU9jBX4TgIhaui0+133SGjWln2OosYS4bgg
6tntAx+uiwclYt8n9UFrZ8KgYk5xGncPCk/kBlA6ew+km/A8TVsRqSKHk6pJAhz2cwa2z694vnjnR6J5cGSkfFVaGcbXlH4PJUptwr+CgEj0pg/r/5eq97ZvhXskIq53
36Eg6yyvMgz55vwasoxtLB7NSyCvrh9hDtZMKSfEp01QdhP3bENU19obsR/j4KiKNuPiF73enmL3njksge7sn0/ZjjfkcQCBjllhE8pYwQaM+Qjz51CQ0y5v5Ghi+EPa
BIj3A69hVRYXj/RJ9VP0MhXIbzzj6MQ49WpA5iK4wWzqWc0805hVRGkxAHJgp1RdpmRWYnSxG2Xib12b1lpSn/fvlN6uTjjnYMJpPEDH6zN/Dsvc6Ule0B5kE3BOi2JS
ejGWAAEr6AMOiHKYhAcirqQu3QxvDBeX3phAFM10Nx8ww6gJn4ytZNrA3AU/W50HR03CcwY+jGA/iuGLUURL0KfcYpd4Pk/KDcMD3qbEd+m2qB4Eazeidzs6wui+WuDV
NtN4Bxig99iVxuKtArz98Gksjy7G93GsmHOKq076yZdJrZLovDPQt1U84dPe53013NocVEpGpge+Akd53TyIWGn7wmtOArYMAGjDOcR0C6e6GQvOFpvp4EsBRG44Pt30
+51h2om/RttbhCupYXftyjvXZYJVcMRTNyve8k38zevahL6fnj1UHvVPr3QkJ+PX1P5rE79buksBPWaXJsufYjP8TSoJ+86rzwCB+OAo7xu8BWP6tOyfVdH8FiWMRkM1
Q2unxBk1az1QSLmPoy2DNDbTeAcYoPfYlcbirQK8/fDzCjwt5TPWmEucPqWw164gTNiD9aiZmz467cc58PT32/jahP+zSjJ8XARY8CAnoZLWX7589iFomjoEf3zgnkpy
U3tjapibmYT3AMmrt5v12/mEPUlDXxmt2hUWIqX6lDMT8iNBbDtpsflDSEBpPhQQuCD+2Hi9tLze9oe3J8+VEqQtlgvq5Hp/YwOX8NE5+nkAcmBid61FsUikVpKpE1wa
jXME+RMUZidKNgjPXTJrUAQQA8AVrXPp/GD6e3nio9dNDpfhUnpDyQGHjbYjPInLnFHWNtQMFQalxoTdZgQjeuFqRmAkfQufeLshHcYd0shOqj+M6B3WcHtiyT7UU+dO
sZoZ5U3MCKJOhTi7e4NnzkHDGQDCZjH/GMV5FnEwqhQZ/8MVhJSRx42Ku4vV01vHu914ZIUIfg47Oxce9Ewe9BCbyMhmkQhuKTkH2sgZDZhNDpfhUnpDyQGHjbYjPInL
MkLhstWIswvfUpQAk2sgZCVP5pETtBukk+VeqIfVmsaW9ZtN+jk9ovYHFEsFgOGkcpAMBUto3AhwrfihGjeHr5BsdZTmQfogQKQmus4E4w0cIw/F2ajU+cPItHCXwTpk
mX45nHVHO/yQzhNCbMBD/i+z958NbHH6oVsD702WecczHap0xxKEuXnGGbb4+9q9i3whGdlH3lODbj1meXIfYVNdpfQe0KGhDnsfLashPTfjT9/Q4dgND8NxGCggNoKR
L7VknNuSIpfpkKWpY2ExlG5UpIzmVMEVPG1z3/hr0+twtXe9a5uHqu11aLr4MGWuR5YB16DIL+BmlIXy1Lr7q6we4EnHfxvNML7PX1ydRv7GxqpF8WSHSq2J1xfBLKbE
duGgTEqUQQ53E9L90TQ/NOjbrGRxqgWZb0Vhcp//NN1wc+IOJ2LnEwZ9PAHXWVvhBu7t2na6PWuxM2wWUc037xUHoPvHajqEh7IDzr1YSmiyuB8sbvAa24hNVMhdshqJ
AcQ0H2TIPMMqiS+t1R7jxMXdf4TIwntBk/bNSN1vcgaQnfaMN2bVXhRKtNZMO4rdhkNb9WyCisb4vNqmmMYyJAuIdzJOIO2Gg1S2FcbXNcjQ+KEtfWUYUiyJGjHmv1IE
aL4Xz+E60hTRKNRm4JyQj41zBPkTFGYnSjYIz10ya1CMwZEnOUHltOvfObuUU6KqUIE0XVn8S/OcDv/mC/HJi2je89rCKOvA4QR0Lvg2i/iUoZwZLywpwYz5/HA1Icgj
2g/5bWH48zghgB0bOZHCq7F+eMVnwGjVxKHZq7BzS6Ry9axGKmRfiP7+gfo+expL4IKUOebvjvk1VPCegfQU7Mhg0wfGDyr6vie6SuwgEGh5ess4VS5XF7cYqIZAdIfz
IqDMAG+fDzWR9vKEDs31+DbgmY0HnC8FWRif7AIEcGWsHuBJx38bzTC+z19cnUb+RDHjoeuWchtQ2BCNkQQOGY+jLutInISXmLBe+u6uxUEO7wwTWc8XMG9a9dIp6sIZ
2lvVbjzk2Y4Lk+1b5pjAbmBzdkPndV6hooo7HAI351V/M6sJXfsSOek2N73b/RJkMwDPDgZ8DXaSg7QSOhjaM1OVXXPgGXpcJMw1T8ZqMc+jZL0eP8NQVsTw9dcl3E/k
GYinHekh+vJrYl4jdf1oauBaeliaO+GoZF9REHtFsszx2laIOuDOShwCfXqPjP3+QgSb1hr5OwlNXbJSZ2/PokonMGI8CtAaI1ajT8NnAUdSMiUl2g7l5KGueGn0jQE1
hDOKTVAOMDhoAYu6xsp471zzsg5NyAtJpOhm36VgeNT5HLIWp4GjNwAbTJCduOAV5xnSHhIBImI/XOeRTrfOrvwK8Uv2deupdm8CKghvT/tTlV1z4Bl6XCTMNU/GajHP
TUglqPak0QnJU9exESK6yUAiwCd+XGI1YqsG094IcFIhtHeiAa+EKdSBV8orvkydyogm0Sa9h4GMq195YwJtiGWVAtS2W7KjfElanIgLLdDx3z0LiY/VB31fsaFDeX6b
jjBQ75PEGCAZy4xAQPPuZ196cpz9eZKcSq5mOlIs7p33Nl+H8uwPqT1Py0N6QI0IlShWgJzQUbnO5j2K35n2mMqIJtEmvYeBjKtfeWMCbYig96O5ZNtO+Zr0ePRhXDnp
zr0PpUFrGHIEKln0/UyEG3E+ofY0AJAlkhAsX0xWlJkB3LcmNT7J2f+rLoeQxTCVyogm0Sa9h4GMq195YwJtiFRXoNxkyWzyNq6Ufwt+dn0WYXG+FnHdTNZPGIst7o5h
E3Z63UzkZrjjV0fozIekWvEzCcJLAM51HsKOUktLISN5ddJbpdIYuTrf6GvoQDhy8Z/HLAP53N1qM78X7/ISNx2yJHGELAtpqaaLNajdegA9bC76X2SPQQDIn9WFXrMx
yogm0Sa9h4GMq195YwJtiKwe4EnHfxvNML7PX1ydRv4PLhI3LJX56Xl0sfwGAF9snkDc3stSTkc77JYJQBH3Uf8AsPGfSsMDaWJaUHl3v7/KiCbRJr2HgYyrX3ljAm2I
SdTHDhM+NZtej3cNgwfItdciGO6KwalbHP/vJWac7OfhFXmAbR6Le3mBWzt5QYgByogm0Sa9h4GMq195YwJtiMiXdhN9pgbLUzqV3TzUOGg2g1TJ4BOgYlSNdToZ/NL2
yogm0Sa9h4GMq195YwJtiLPqzge+g22Bp+dJaQJvBsDKiCbRJr2HgYyrX3ljAm2I4WpGYCR9C594uyEdxh3SyOPfXvr60kG9g3gujG0ZDR4CtoIbqs6JW6jRcAATcEwe
tPY34MKG65g+dxI7PnG4vz5idZsBs1JEZM2VTzzFBKo8qpVohIxznQkr7UWhXUMBWxl1AC108omuYnUm2r/X74vv+0sdQ9IRSSIe0MBUl3vKiCbRJr2HgYyrX3ljAm2I
ObbfZ/whuBKQLD5mX9N6UrQxJvsDNf4yIksSLkieQUpc87IOTcgLSaToZt+lYHjUyogm0Sa9h4GMq195YwJtiCKgzABvnw81kfbyhA7N9fg24JmNB5wvBVkYn+wCBHBl
yogm0Sa9h4GMq195YwJtiLPqzge+g22Bp+dJaQJvBsDxMwnCSwDOdR7CjlJLSyEjeXXSW6XSGLk63+hr6EA4chXFdsdoz94eHkH/bkJZeUeisaUBY202fRxGcSntmVeO
m7OUpyqr9qjffPe27Ox6ApoiPd+tizCzzWWfZtpSw0ZgRy/IQGhzpVcDZVHlfQdX8p2FBN7SzPVTGIYvNT+7Zkefba1b0fX28iqjSHn31up/VeZZ4oy4xZ+DvK5CEUNk
O5FWiVFkP9mq3MfFH3v2FodROXE3bkqSSQcwHHFpAV2JecimXmtXcDsFbPa1BRHIAQSfPquL4q7AjObfAaJ5geEVeYBtHot7eYFbO3lBiAGsHuBJx38bzTC+z19cnUb+
Dy4SNyyV+el5dLH8BgBfbJ5A3N7LUk5HO+yWCUAR91HIl3YTfaYGy1M6ld081DhoOBmPcbWoYUA+M9Deaq60O3ecfunbe8x87cdkgnSRS3cNPRKdgbR/ub6Mr9AIDgFw
xUndi6LOcsGgBn8zknXvH+Jw5d4OPhfMMsw//rht4WfUDnsrukdBnXHlvHZeCYnFcpAMBUto3AhwrfihGjeHr2wL8v9zeG3Sx107Q3bLQxHDX/4hN5+/+rL8BZzVIsMP
Fol2CBe0GJJz/O7IyvmYew7gueiqxg2o7/P9tfOe66wy0l2PWZYWgSam3S4VG2KcY0Ld4Ou2cLddGwXnv5hcbFr3r6nD46n0gkfFSgEEDRdPIWfEEsIV2qEHc8zdFqsi
FXnih4BybSSj5IapNULV7JCXtHUbvcnUrHQDnnoZso7qK7tylQFb5UcljfBRZhjOCiwHhy3ClQmFIDmNbu+0kpT+vrFNLbK3CsVZw3M20qeb2BNh55TQk+b8gwIF7NFp
pYHf57NXehryHozM8LUjnqkZMm8Zx0grlM2t8h+ylFyKSzZf91eZ5LQDWy4KYC8tU6EIPO1I/3Od2gYUIGePln0TtHxwqJJ6OEwPjktvxqfl1YhB4W7gMIslNVqN9TC7
BEPxcLiNr2uGwvhboSJH74IMRbYL1gxRqR5RmsiwH73SU+4EHT1TApR5CNYAOSU7BEPxcLiNr2uGwvhboSJH7+eZripDF+Zk+xqGaktbPnMqyjdVeKWZ7C5NaCpXSMrA
nJ/ke6EXREq9YL0GI/SkXFLZv6NSScIIX+x98us3Ye0YoyrtvDpzJioFIs/d+WVEPMHzd24u0LQ0OneCQJ9boU7DNxVzvl4rhBu+45LF/1vSC77SyJmCm6nUDYygl8Fl
BOaQB43hlta6j7oPiu1Csb1kVCqlYRYZC07/5l5IFE4gafMhFhuHbn2i+Reiu1msJyIJ/TwHcVIxkrGwbrBPk1gF9GkqvI3T532KH4N1qB2vRCaMKfb8q26yR6NXzAUf
r2Q87+JnL2lDCd4mKOi/6kgEQvtW59AGGvhXnnwdHvdToQg87Uj/c53aBhQgZ4+WIBMBBalGK6Bz8BpNwVKVrWSNvujCRsLrRe9Ukc5bPJQg6Pxq/SSL1oHbgT8lYtF2
x0ouf1SR9TYwKuJDe1GDI36YZkr2qoKL/GiQfrEN1/2IO48/gSOzg+NSkL+SrZX3SiBrMzsvSgjnjzp5z6xQ0YsnZXY+8KIQYQ74qqtSm1DdPtSTGvF4S1QdLWuImwzW
ov7ywEBicN5gAXl0VWOyEq1S7h5BB8E2PuIS/H0pfsteNFw3lh9He5DWASrbVtcg/YBi42zEShgO8IGmJ1BTxyUy64jEo8O8cOgwqXHvueUp/Bf6z6E9UNbXlENtP1K/
cKla5H128CedsPji2kaZ19iruEB4IQY6bO6AXPQH2jjVwn65RQO5VHjyh9xFWRs7bCAFk2IBxHCteELqy5P2ViUy64jEo8O8cOgwqXHvueVLkj+ArQkgfNAbzqsu702p
QIjypUprfEh+A7CPGeowymVe2hVeNUwX+QYHGSDcWII1MkXu9cRuAjREJPqMxBrhOAXLunYBn2I7uEwmBo/MQGVe2hVeNUwX+QYHGSDcWIKS3TNyhPd2zXV5rP+WSrjj
sL+l5ixmlP3W5K+q2vbiZyUy64jEo8O8cOgwqXHvueW+u+4qyEAGAUUmUx2HyUR6cxryEcozxNSLhS3YDpFWNiUy64jEo8O8cOgwqXHvueWjE7+JbUAV83FXqx6D5973
c/OShjgnYDBnHLjISR2qkbJI8RgYNBJ9F+hstSBGRYfKNKFNM9YQc/P0eTKPA/qiZ0r4HdZ2IY77KHESvOjAKyUy64jEo8O8cOgwqXHvueWlIVbAVE4fjZnAvopQwdXj
ZOfDb0YOZlyjO4u7mVZnNoIn1rVNId4cRcwiJViwTj3uQM7gEkOpnCjBhCd7+1pb3vc9aqxMGeFpaENZyuJ9gJ9wyi1FWXdUaWnJftte/Px4QhPWcu5MyZmcX0Z+PNUj
LmKRiI2lIu7X97POMWrj6/tWYGg4OfrobgD+3kq88spQ4UnBkDIrATBm7se0jqV8+T2w9EQ2sWbu/l5M4S56BMSx+FpngQ4bI5T4gOepG9ZQ4UnBkDIrATBm7se0jqV8
JbwzNFKQwakGbPy1FcgitwLixi5rjTThTaKqfzXNbxtz85KGOCdgMGccuMhJHaqRxD4dj6qtCVf/oHiMMOjruFV43u97fBaDFkgtr3ceufVQ4UnBkDIrATBm7se0jqV8
KTEwZGDXGFJDW8GRGWNy+b+/NGviR0ungZUBxMhuRSXEmBPSk0KCZ5KTVBLjAZeB+DDMf3bInXJj3pmztFbtBE6eya3tApqmc6empqiZ71nEmBPSk0KCZ5KTVBLjAZeB
Ev+RJsAtmKZqF8q0/Hj9hY1m/MbiPS9+NJcu4NXFg4NQ4UnBkDIrATBm7se0jqV8GJCKhVWPqWAsY4KpVwW9qITeS4VNEKhX81h2uIKsKxlQ4UnBkDIrATBm7se0jqV8
0OZX6XWc4jbzoVY649zGt6BE/pXrjj5JoRQsERpjziQQiSzkvh5Gw/r3o4FAFGHBr0QmjCn2/KtuskejV8wFH+JtMnxwH3oIdQAVABOREcVQ4UnBkDIrATBm7se0jqV8
IsvDEyu1b2gMeluIeSJ/ZgCvYVRPtaLr46WoLDubj5BQ4UnBkDIrATBm7se0jqV8HE6t1dTGrSYngr6zsHvZiyJ0hjXmnoGv9PN17zDkLlRYBfRpKryN0+d9ih+Ddagd
3Sr0kZ2Lz1V/Ezom5fjrHMrfzp2LFqEYzIW14ZHqeXXkxMfAI81yez9oxFeMNsTe/xz3L3vPNgR0z6hWJbn2p+IePStPGhnptG5vwBOv6+aLRbcOFMdBjo4+1C4yAMIz
49ikr2KDHmwGGOooje69z0Hnq6h44UPQqpzxmtQXUcJsXu6ZenGomReKxh8vChIhrJDYklqdNovF9fqXjIsTI/BkX87ESeMxd6hISZdNcgksZYcnCE9FryF0E7+G/DCa
7GP3t4RQWWcTirZx14DSOhbx81m4gmQsvainJfMzdb9Y9fjOl+G7Cvd6ePZa8sba732R7rBpF2oRxxZvbB5lheS213FRIdUGxeL83xJYGCg0PSJgqmCg7zpgGkQAwuHB
U89LEFx9zFW7Vd3Gc9B5SjYOSBfR1G58qYYL7WjxkyDMrD3VlyF325zE7mZMXEcdC1W+Lxy1OUG9YbhV5ywzxMUIFyzEci/VfmUShRWDyVJmDG3fPGIjZVYVA638gihu
xgZGBM50G5/+MNGcv/PF8artKshpCMBJEDAbkW/fErcYjXC4aYWsPE6qRbEm3Gfj+Gz1HcG3zSZn7HE59S8LgII5K7SyYQYLpfg/Hd3xhl3XFCk422daw2+KPHly8V3A
VE3AeUKtXQfhrcvbmFFe6dau1C6kk6k6eSXKQUxfax+xs+K8g+pNR1vHRMWbL3it7D1ExQPARZIy6RWbMufF2wbc0Iotb+xflGPgJ4f0CmFkEeA2/1Y8wxBjK7rjNjcE
Nz3jyI6iXf2J5ATDX/TDJs5WMUpLSe9xLW1NqApn6EjAtFotYkDbx3xv1aJsQTkVgRHnZKH7nuOp2D7SQ1hZ9lvq1fn8bIrNgyG9wn1Bobyii6bAVrvDv2smY3SbaEo1
xAkQDWzjmrGZQt2MtkB91kAnneZCrC9Il1Y6+yxSFc0jPlTJc+aE7PSzruqztFxmN2h9WQittkAopxPNno8HOdcUKTjbZ1rDb4o8eXLxXcB0nE0EmJDkJ1yYTPE7Fz5F
P9qrET6eF7PH4vosV2V1J7u/+n7LzCKhr356aUQsccnM/Y5xq5tAsxgPIE6tYk7ZBtzQii1v7F+UY+Anh/QKYYjSDfNFbBswyPOJaQXBO/D1xyL/L+LzkXkAa3e8AmED
XCyu67aNY9O+DErNaa7a8sSkwuVTce8aLy8SBlpHyT6BEedkofue46nYPtJDWFn2/vI0VgzY3z7UYXleyTYTl6KLpsBWu8O/ayZjdJtoSjVriIjh+mCl5figm9YiPZrF
8TbFWB1pBPa+xcyqYYdt8SM+VMlz5oTs9LOu6rO0XGY7qvivTe1qrfMvkPampaG2Vjzr7BAU0GGdcCSG4e23LEOtWst/mRAcYNpS2XEphI31UtifBtCMuEjehYrbqU7o
H4W2ehoEisrLclb1VCRTg+YOnEiXFTO3MDOWzZI1Y7oV9FjiFpz9o0SBuYUgxg1KF4R6tRg6jPYjY3L6VPitcRtf7jr0OdLnQHwI93DMuqJM44gFukoAmWARZ0SpHBmf
rzCfvwjuOaUTNkwrom1/KDNxLvdlmZhVf7X4IK/Ap41PN5EPLPE61aket6PlM3cypzyBha9Lrjka9ESbPeTdymegp3bgvBpqnSFO6kf/+YKSrmg8mVa6IdJhjnkljAI+
FfRY4hac/aNEgbmFIMYNSvvc8mmXlSGKTD/QaTGyUq8jgQ6HEC8bhNaXki993q7Ac5cn9INVj8u29SDQMGLiivNwwVRLd7ILu0PZFbYxwuDXFCk422daw2+KPHly8V3A
zilpdbtv/nX0MSRs2ZKjtQ2DbJ0l02GOUtwY1dQU5OWLlceQaWYGcyScpdhrNQH7Dx7EmTZqu/JlLjaPUFAuXtOk4zd0yqKQYeOvpsCbqq3fWUcJeQCvmE8P8d7FkTzw
zh5pjVsFI6A6TyZWDBvCMW7etCytxCaFMg62Ga6lE2ARIrqk+FLQa0uFF6+W79XsM78g/OAaHKot6hIuCzn2ObsegXPxBRIA62f/p/ZDwL4V9FjiFpz9o0SBuYUgxg1K
MLbNTd2VOcrPl7z3Ank3nFWt7wIspZULibWlllXpXJFzlyf0g1WPy7b1INAwYuKKOxFnxexJdNZmiZ+Rg1UquNcUKTjbZ1rDb4o8eXLxXcDAVtliz7Z20OH0UBy/NIp/
V762aYjw5jkifLZTPkeFF2yfK0/yMkGkY9Q91jhya8Rdqns1a0fCdM8soSzW8/9+/3vQwyp8Mit6vANbO1OFpll4ZiCUCNVVJLPnc9OZShwp1c7freRwu2pAc5pIP/Yz
/fBnZ5a31hh4nXdf4SNfAp8FmiTCF90lCl9I+aAv4YHBQWsbBniWTj5lOnWJrVvtaYwMlnn4Fq+1WNGGpNo7L6tePDCDaDtIkcAHmDROCHXN2zbtICS7LPpyY3GIS8JX
eXrLOFUuVxe3GKiGQHSH85TPSxQ5OV3pn3j0I3adBYhR8ebmtjMgenXCYNeUdNzcZu4WUmgiWKMkx5Nd9Uelv5+BrfPvF+1dkWEiEN3tiGdmvsMPFrUvd6JTQPKo+Mx6
GdC30oHJVEbSL7chcEC7vqBRWeb+JVTZQoOUd1k1d/g4eZm8yFiEcLAQ8NFm8BmYIBt6IBH7qcXdWaCiQbbWZMUkj8MsG9ulZlhBqW2M4f9wmlKnPLF3x5wKOoPcxqug
ZiyjotBm5QCO1JGNcEdgwQcn2SgSWc+9Pro93WIZq13m7+uOVMv97PbQnMtxCCa0qXF3M0vq+PfNImOushw95hV54oeAcm0ko+SGqTVC1exDzirZU0JeskKO1PiDXSDI
I+mWmaw/F+bjlRyhZkOvd5Ul2fJT8Ot7wRMN2b+G/5vS6bRRRmDoLSNPTmtV3AIkm9gTYeeU0JPm/IMCBezRaYMr+6OtXhHpRmnvFSU6+lA5l5GcmEMMifc29x0yXyC6
kSlfj0I/haoFEuyQABotJDhxF6Q1GJ7xHytgvc9wEp/K4Gz8FFMSXpZIKQAOGQzTOQn+z27saTsf5/vBGJysxurvyGXlkWCRloqOqsigPDeb2BNh55TQk+b8gwIF7NFp
qDOegbI6lz6a9UQVm6UFjci1WUDf+xFB749ou/IJAnOXXZqNtMf5cN4NXnb45vtI7hqW1Fo1IQj1fuPf3ltehRCJLOS+HkbD+vejgUAUYcGFULktOHFo2ar+AtXZRvVI
3GFHBTUo+1vg1ehYuNUeroYXWjyCuRIfZ4ijWpUN0DwauInJ16QAM2/BPgY0VF7Y/b0zOe+ZL7ZewMPU396KESFBkWsDkaaZm6McbN4NPQ7U4w9I1JQxCOa2v/iXABWP
WAX0aSq8jdPnfYofg3WoHd0q9JGdi89VfxM6JuX46xzK386dixahGMyFteGR6nl15MTHwCPNcns/aMRXjDbE3j6SUuCXwPf5QbIGZMc3P99kjb7owkbC60XvVJHOWzyU
IkPziNZ4ePQB/VPrKuWbZHSbgQQb2ZUnXt1YTk4A5n/kA9b/zIxD15cW9ijNhMwCPiNM1j5TB1kmTEVmEWdtOJ/Cp5FViS0iU+6DKldMfx3nV9EDXy8EFFW0U2D2680B
LspfWJDhrF3VGYlPzzcnEiFI9tBXcYOSjEk5I3rXDacqwTonvIdvSr834KHjIgrGsXvSfcGxEeZpp4gHWh2A1XjnQhcUW7b5xLlEBxHdwRANBz4LtvI1P0SdahHCnfCP
JTjqbQbhAptCFNFOjdWyVwstoK8OZtkuBZ4yStVXq0xajuKHzJJ9mpXwgaFonJkr5rHBiJYRof3fl6+emPRllOPYpK9igx5sBhjqKI3uvc+HPjir6VdAi1Vd2Vy1GdA3
TnEZGA4GgFoa91H8KHEO4bSi42CibOM+/jEPGNo3WyMXaxjxWybuGefm00d0qcKyPTb4bmBcd5lMtSNG36CzfPrTwf3ewIT8hWElR01ZUAV+UwLkSYsavBbUe5lmaUo2
ZupDIWHg8qsDBhhhqkznQHBr0NApGRY66Klh4NjIjl8qQdNgtnd4VWBHoVyrxvys3at6LdNMRL3OTachB/s8DLeLaJ2f7j7IBdYIP23B/Kt98Id0+Nex7IB/e/C5Fhei
vt2KgEQN0zYOX1IiijFVDXGlGl0F8x7441Pn2DqBrdKxe9J9wbER5mmniAdaHYDVn3mNSOeY3xlMG3KII1hAgilZK4Jfph0C6WJsD4NGaZBCHhZ7dUzUxGofbZ7MXoNa
jRWTzF6Ip0stanfEAkzc8ACpsNM0OVAqXkp5+9vj0cIWWb2CEEmkO/Q2KLdnMNCtZ0ph5iysJKER11Eget6uRYoO6e/mTER4Qs76ZPXkki70cbwd+s7OvEF3Ro4Uf2Eu
BPP1fAEh50HNiLoRBT7zOnoTAd+7M/7UGvSZIT602/tSNXj4ia2amWigTr32225DTysBw9sG4hMaK4+661meXswH71xp2I6eRNDSVOhy8Xov6aKppCV9iZTYon59Xa4V
fIkcyz9+nLWvFsmr3t56UZDdT2rcUC5+gEQ/BhhH+/U/1N1V0fd1Fyfy/cK5RuLoyogm0Sa9h4GMq195YwJtiGQN/riwlph8nCDIXXAoorcCIxw2UaC06Ign2B1mlC4g
tjLRAQXrMfLV1ASaL50f2b7dioBEDdM2Dl9SIooxVQ0ezTvGU26F/3GAkxHFI6CHKVkrgl+mHQLpYmwPg0ZpkEm4qQffziqpIkFJouL/DVNtnnJtAJm1sfOl4QlYSufN
Qtfv9p1+mTuhRdzIqynRyTZnQ9rNyRUW53gT22xI4B3KiCbRJr2HgYyrX3ljAm2I7KvnkkGEXOxhB8kOFUr2abEX1WsGHTf/DURp7xfsdwWx81MSaJ6sx1W1pCuOfhKK
UpEJcA+JoTc5gSn25PctGEm0d7dBa2K+n+Gy8LWFKfZtSkhKIH6rfAqIHCbZhDvcwnhpVTvwwoJr/ftGExDiE8h880isrUdmbYb/ZCtBQ0WShFEPum5NWjpCgqaDqsAB
HbO63Zb4PHaczHaBEn9NWE9N/krgtaxCbaVjz7Z8jyH0AJXb5rnqcj9LlGEc+uCp+bGxoRkZxImnbdGBFOdmwaOKch29OF80/sWzDERdMUerS0svqVgyXYqWDun4Tq7D
p6YSUcJytOo+nkdEgSdrjLrNB/VdRqMC9ZY1+vDx57zC+vxH0+VhWrPKE9/u+wgjXos8P2OT+IqvWafeeAmPt/D7mQpDWBMYL8h1Z+rqBh2liB2jMIT+dmoADlfzDfsv
VqTbuBt80yfhLiqlJEkKBk2Dfl+hqVJb6ihdtbRaP+6TjeAWkRgd2U+EK9P3ldJJiJ5UPYnaHikW9FcnVYws62oxCCOpfw/zIEaR+oa0DvTyDGAQj4lYc5ksE5ypsty+
5kTHaNKTUB80BmhsHE6nDWvTc9Z2Q7TTu0dfuaEwHY07l6+MNYRkJGkOII0k61hvAXhTxLNQm9Rm0/aVcgvbe4+dQ+MRJTY2Fo478hgxqyCddS7m0N6MIUjcWdyOeVvp
zVPPtjNeQQ+24mehRxwFF4cGywlmV0fqsc0S/ctaloI6qFj6IBiq18B5KPdM7cC+Xtz2fFacxULB5FejHsD+IdZ2PS8H36DETzePr5Q/YLkamnW3/x4T2hmCTlSFI3qc
D0lUwusrKXOYNowDYRKDK2fF2A1gpy6tIugCDgN0ssLfRQTmaMreGV4ST4qlKN5NXaIwOGargKESTZnVqEqxyaVooKDyOMF9v6ksORVTaswIZtzkGnxTkyb8pO4j2HjL
tv45FULL08z224yvIMq6g1hJj/sJC4BD7fzjlccuoW1kFboHxZsy18HK4jR7W0JAVfdxcVqW+wQFmzN0KydupcqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFz
qhmo6irnW+WPKa7tFrq3ISjyvbvoG8QIcmOuj8u6Q1rZa+2DlD3zI/oLS4zu8ubGyogm0Sa9h4GMq195YwJtiNL2fwuQ+LsVfIRkdOsgMXPa5MdcUVse4DAV/AcLmKtQ
KPK9u+gbxAhyY66Py7pDWle8cPoxIYYnX6OxgsY8+vuD4c43ulkHlsjyVirTosgUSeor+1VsbbG5l68CKHhk0hUILneXtFO+h0anLQTjycMe07czZ2duKjmUJjU4wmLj
BoMiHPw5GySYp51IAbs4wcqIJtEmvYeBjKtfeWMCbYi1ae5gGLv4VOyVHTA5IhxdyAwuogtAtHOIvSnNzuZuk/7opcw7Vcxv79sGHTNEnQVCIf7qwLt9U+/9lG2X0qvj
FQQthzNwbX9vD98ItFSrgMXPEU7ujlO1s3cVlWjqZDzfAffdedpGKq1rXSGXjvLas9onqZcWsUjN8gH4tbeOfmZPUIaY8nnHEEtsz52et5d87h4Xxj9xw7e8FD53Csz3
bj3Ko4+CjH8yg9uuGxmZnU9AHUqNPiKMXd6TmqYHnDGQCER9dmVVn/fLq6032MyJAPnhKkMwlqfLjKsd1zmACvbUemk62T8t89BbVyUm2oK2y+yTlxP0KLpih3W3hj8E
yogm0Sa9h4GMq195YwJtiDpnAWVVHivKDTBw8yw4csFpL5KcJexzrz2RNIP0AFoTZTZ7Dojf1+m6i7iMb9AEQRaRvOFrEKNjNpVvAi+x3SGD4c43ulkHlsjyVirTosgU
Seor+1VsbbG5l68CKHhk0j71HTn14m81fQy/PIbQNkR6ijmp7TPsHk8rdG838NL6TazntDzpZp7xB8xtw7gHPt4ER6ENG7m0FDD1bgBFTDrNXtLtfDARzwmVP2fLjDqL
zryH3oMad/wXhUl6fYM5FICjv0vYGEGhB3hfzRYrxHU4PsN2kBr0hFOZn69EBTTQ2188g/eDKemq5iGUgrpAe4tlG5Ew0kEi1HUSNFn6amS4qrQZDcwWujDcuwR+FUoV
a9S2rnBy+HEubf1NXt11wIxNIC68cUokBxjrq7n/flv2Ep5WkTgLnEHmzE0Yd6l7+h1jrovmtBsYyOo9hiv1/I+GvTsfC+mBm8giDvrxYlfuALI4I05GD1cOH1rMKygR
PJ5sxQVu1tb5ddc2mJ2qvrzXHGp/aXGIqje3skA36sEmUzt2K3pRXR4drv4i682ouG14LMm1ivUYANfmj8mVVuDPZuO9djkl35LByXUAg9KRUpGdPuXkKkjvDp9Bmvu1
dnb1zBo8FV4wlIP6eaSeF7QMf+xXJNh0r69qpCM7xNHG1IRyJF/DfHPl9i9ZwjTZgq8zCNh4hJeF3T1jKWc9AT5hWv1ogt/zGScYLvuLS5aKDunv5kxEeELO+mT15JIu
W4pii8num5x4vZ7JotkJaOLQR+86kQif0DmF+si+6kas6L2sf5u6X6GaNQHXejs8xaPyYKAVa84LaiSthv9Q5+MEcrEsVWSF1K7ozuyXe5KHuVsaZSVNnxweswj5EDyh
gq8zCNh4hJeF3T1jKWc9AcBRuAXvBG8a+ZjEAEBl6wJjpO7v5mQCn74hlmUTBoqlQfX3OaMwu356fr0/Bmj9wrg8awjRmRz5VTXBYRad8eEWwss068DaOOclbgEiVuXm
AJ05o1ZaGNPXdDDIyLFFmRRBb0BWI4fB0MQx7/9zmRkoPofivpn3/NExapRGXajCuPAub5ggWSQZ+Ldv1bJqp2R4Cnft4DY3nj+YJWUbUXUq//uF0mxB3QGDBNMDg48C
7AtyzQzNvLETWC95TLdXIFMU3d49UE+tU6huyAywZrWHpb50lKihrcxb3SCBDp9PP53HUuDJ4bdvyZ02xdLaY1SBnytu5ae9yNhkaGU5NjnmqukwF0HsJMaCiKrc9lpt
gNow8BUcVzC/7DBDqqMvrApVp0gQBqfnlC6pJDzQI+T2mLCBn37+TfAPKuNGtXzUaO7IDr3YJQXD5Qnr4jBj9GY2iS3QpWNqfIhcyxyjZjSNWDMer1yAkn8TEqg6hPf3
aTYBztem0/YbrNkYRTzQdvY3185GL0I3XIg2IhFYmB2c6qZVVHYMdhqGUZMgbba9rW5WA5LRXv7d3ACExS+8v76yWYVHC0c0nIqh8riQkhQCW+8i7BfcawwsS1BEeb8R
gb+5zShYP6VilZg1OxXEKVi4NIhOr01eY8uwLbUsc+xcPDiIKBEeOv2WYWiQ2fgZewbiPTO+zy/tubmdEWu8JRg5IZJ8HZ3UQYtOossRm3cjj/neUe/bBx8rg6ahtwtB
g7tiIrG4XZ/cqflC4/3S+pXIFCaSU7CQrUjmBBC23PqcNXfx2Bi4l9MlW8AQ5yliXK/rLMVlIDM3U4Pvjrky3dmJD+AQIRwe8okxIkLiW6r32sYuM1PLz9SoqFe7w/mn
rXaKXeuPBvWiQVxKL/quFQWbT75HUmkiie3T3SU7z1oVFbt9H2hyClrX1+3YNGmYxIYti9IDg7ZIOPQ8g91opgl7ofFsB/N+DadQOj7dWmSBS71Oe5OQfc5BtJr/riGf
aj9dH6YYo0nmV2Tka9lcJL3lPZ/wt4w3M6U3K+NrcGCbvEV5I45uyE6dOdJ/KR3WWtj7J7F7POZfLAfqZ4n8E9oDyZLjE7k4I0bgXH+0ZWT85dW/LbOMHOJPp1wRrNaf
T6yH5qngl2ynyShFkobDjr2V5GQPady7FuNGtCvN36FZAR/TGMCghkpkg3w713SPExJ3jSV3XNjLQuWy650PQd7m/FxGlbfHbkAuA7dWXnZJJi7MCuK/LTRX0smybEi6
6getE2U5ItaCH/twYylcgruxjFWFFk8yj70zmdQbFNC9R+Gi5ZI2bKSVv3bsiS23TMOhBksEz9x6pscMwVmFywhEeoVSZ7s8iJC9OfafE2W34zoXHWNcj0CXXcb7rwAO
NCIjw8qDU1qpmu3HN7hO6NZ2PS8H36DETzePr5Q/YLkFoQKVvhZ9krM4qR8IyaGueTLNMbIKKCScOjn4/1Gge+3I3DKhEz7Atndj2Yj9C+YpZ7ChROSwiL78t8sl7yp/
r2tgvDLBSHyiDGo3Aj4qqSlnsKFE5LCIvvy3yyXvKn+DYXFAxXG7kadVLLDjKrkR7ZAtWbCeVEI6yCqugXP3zTujrlKhY5r/R7T2LVWxBxgC6FGgqx8aVMD0PwwSxtlV
Z6YqO7UOX2cbWnLGVDUR2uEVeYBtHot7eYFbO3lBiAFCHhZ7dUzUxGofbZ7MXoNaJ/0ueG227rIu9XCWdAFy60m7iOJeuID6+2KFSAB/Sn1XLq8Ruf82c8pYOXTIR4ZV
jCaIAgj/2+MSP47yseogwQ1v3YqWKquzTTF1YIQa0jTxUEsXz8GyUTJuzajC9ZqX94DAdFcUKR5ko2XPz7Vl1MVg+tkPJ/Jj+QoUubfM05vgFdd98i1+l6eWkLsbMpto
Q9uo3RAOejD7yPkFrI1wZbXlX6svF3DYsQEEN1ggMim+m3wD0MOHDZU59P8w7CCMbBa2FaNyCNYpm+HzpgD9E4TRDm7o2Gd/ZDO1myC6dAF1sE9aGu5s+kRqZbmS2PG0
cFmlQDDBWjsRv1FCpLwpepJxzFcoud1Eh/7Bg6Z4A6SeG/LFSWRnMjuZ+QLJd4m4sEqGr5FwNzh2VRv7OHmwm3dy2jw6Pl/Bi3DAGs5oPwApmf0avsavBgp3jPzMs4u0
4RV5gG0ei3t5gVs7eUGIAUm4qQffziqpIkFJouL/DVOm4Ee3tvDGZ8SkLba4MttwuPG4eal7Ynz3ykCY+NSSPMcKUCRLM5Y7PAJEFjnvp6IiQv6Rz1mONcz17PVpYHnH
Ew9oshRs547tkMtiASEcG0FHGb9UMjrcjLFgEw1YFaPIkDj7gTtXaFg1VY1UHVl1pg/OezUlbP7OUEejrpY0+9c61JSKTpHplbGlHYHxJUbgFdd98i1+l6eWkLsbMpto
jtdUvTN70oHEYeHOghu1I0YpqUtK8mXa8rkZHkSdQF+krxtLZAM3QEuDuTIbUWuuWorFZiZ2n3xSQOOaTQ1IECj6uxnIM9PTrWiAduI+c35HwDTaE+MBSftK5YnTAqIk
a45AQE+CvRbtELf1zPnpoj5SUsdmjor6yYIb6/mMt1LK77RB6IEtqVOQ2ENBHstx7Ce6aYeKgRTWKnhfmGV5OCn8F/rPoT1Q1teUQ20/Ur/M7qa0K6PxkmMf0pFbMXyl
FrqkgyE0thwEU7ljKuYFI1EKQ2C6zGNvO91hguLYTDZ33Q8G/cQi467J2wCaIN5Vd3ZVX5LDasvXFGwOrgHeY3SbgQQb2ZUnXt1YTk4A5n/UIbfQtzPqFmTT1d+Jk2i/
U5sfrIsuBQu+vYP36m19UEVE9uTbVGDsh4qYVke1I0fdRN0gfdVEmA1cUBAYh0rrNWEX6pm2zsdmNMp2IBhXlMhhg4+YTPavQWiDAEBPBeh8ffPCXAY21wyL6/CGuG9u
2RSRGFSm7XHFhiZdlmAk7UJG+OngebaSaIxfHeOL06JnSvgd1nYhjvsocRK86MArDibjyXXLJX4mCEcgW5cauc193Duco8wSO9fmjj6TBW3dKzQBErxYtdnAlT815O7b
gEdaVG2oxnQ/fXlfSoGAgi5ikYiNpSLu1/ezzjFq4+vvbH3SRvaq8LRC+/RDbqV1tkmnGZgjgN8ZN+0nlA3yoxzM5G4xy4L7NQMPm05xoSn6RjHZO4gRXwninCwMLL9+
1DUGssDjEHO7791mUJRw8pJ1XxYpJ4CBzJILILhMHsefE+scFMOBtc8Kxbw51WtbRMe0g7shdEuSAHNcBohXCTfb6VtoXezUgm7FNb0ocv3bhlD6eouYkncO1oohou0A
7PM6cbzV9ZpRfb72bmTG91HXundYlUcuJniCY0XVo7GPZrCjTIO+Q+vW6P+V9mJqRfZg8CBEIReZWrJYrOQ5Nh5nBMwLT+sElcLlAqzq83A033OyMRulc2gpAs2u8Wff
Io4P6aFwhzCJgMRrrMrlzE4BEKgUQI5gIgXstdOH/Xu3i2idn+4+yAXWCD9twfyr4tcfc/udVo5gLmqj7aw4QZgTfLqRlhv7pRWcHmpXldKMdBDhU1qjcJLuoyp/Ze7T
QHCcAaHBPpcQobJ1YVjGtUTHtIO7IXRLkgBzXAaIVwkySkRyCpO6CkcyRwDInLUiR2xPEdIx7xRpEQD2z8jxgUx9mZPMZWfpLHxFvDCF4z6EwLxtAVNF2aOSOxZghgIF
wnhpVTvwwoJr/ftGExDiE/EZVOJ4H7+vP+C0rBZ0M4FnPTDNm/Sc1WuCMa/B7L/Sheb4fbLXm7pnYjyiQDO++7kx8KY4+d1ecv07IoviiAU5a39oVwlTdcxCW7tiDXVM
C8SHn31cRjbYodJoLWhJT5nn8WXWWA2uFvyGVNNA1yjwzwxozZevVGkI++hh/8RkJO3F6PUnvj9mTd+cIUk1kEa6BDNp387rS3IzNKsmJYDDmg45/lMHZThx6FipI7bJ
rZY+XdSkH4lY6omSSWNTVxajEZ1wlVxkALJsvqo766SEwLxtAVNF2aOSOxZghgIFwnhpVTvwwoJr/ftGExDiEzSoCf4wpHGL12JLXt4cQ0WVgp+hRyZsupQWTnnuVn+5
Hy6LiIlaBViKDXy78DHZx7M3Z3nRmcXcKFZIxApeNQlRvB5ecLt9k/oizvFdXTgL4DVR62C6aIB2Klc/IePDTeTr+h2VemAAaUqy298zl6Xf0qnNwTT5xGF37O8s7/7F
jRo1myTLJs6BmvIXX0B2skdsTxHSMe8UaREA9s/I8YFE1lmjDeY5j2MG3BKswRY+yogm0Sa9h4GMq195YwJtiBjB/17G3jSOvDLp+PpSUmpUTxnPCBynjukeCF77ZUzA
7Tp2hS4dNwQ2GubOqiYZZEuQ8RRVJEWgtkZpsZ0j0/drqrXShoY9PlyegI72ZgXQjK98+R3LyMBhgr3XT7REGxrfR8cFxlUGUVS8TOr+yU3tyIf3MQQW6bxIYS+eKsCT
C0Rf00a7gbzqg9A+2pCBUdXKu7Bm11usOE5OujffFdvjDoNvvhHsWta6JSP/7f449K9m2o2mtniMesGXSOhu/JRu+xjKqlMYQevXpyjngq/GQlUxQUms+pUUCLmQDBzh
3/928e1eQpmI1P+2CIc/IXjFf+6q3fiC/j3/JD86jmpKf2fkFZw7PgW5FtXKkFSwxSQUpb6+KyXrYWmgg5yMQyVHm68s+6pi7AGSf+6ef5VXirV1hQq1AItTPMScpjHO
EqpQsd3HjKJ7YxQJoH42AaiBJDh9urUm93XofNC7DVB4pPoIXKEYSxE//JxcrkFSxbyca4QrTbIiJhDC4CF+ne/z4Mlo6lgjt6oA0jUF4Aaq9y4NBELKDp0Gjz1bEnvQ
p+UTsu7q8/F/FDvxFQk4wpadMmv/099LaOxoggBn3dVD7DTU4kl8qHU3ktAHrrzYy9SD+Wl49fn9WCFuu1TDcwY6PpwFcdIKYIj7MOfNTT1nxdgNYKcurSLoAg4DdLLC
79OjoE3ucIYUWnLbQ4MPOapmB/VKu7S+Ay0kh6oSkxsxPKtuB0lY6EmWUnaLm+0xvXOIkLaREBiqVAf/c0Nxxeqrlszh+AtsiIgJ1mMGVqzHKq3eny696++ufolCitf/
OGbJ1XICG4zI5ED1RbqwjrkCTnx/l09QsazP4cQQMJ9+cLv2Nb5BG8StQN7DW+p+8N1aPxmevwymdDSlfwHvUKZP1CH411txXaF3oi6vqSykzClCGoXbWtM20TbCxsiA
Zc4H2GOZ4qx/SfTSBsBxyvNVdTMPLuDTII6axeGqbd/i1x9z+51WjmAuaqPtrDhBgnlNMsgemfd6gFC6BLZA1fKfhkovNsB+U1LMeN3VvCMdbxdAYTi7fuWGND7U1ypy
pD0FvraFEh2Z0G2VL646M0OhpoAUHo5k32giekmsPubq/+ZBy/2Ryb+OXc19CkqsubHZYn3PWNMGF8fqH43KCk1lT1sH9XqSl6EGYXUTJoIB13kdxgu44M9U0jvoW6xr
LCe7Yunj7+nqNkxwXdOB0/Jb2M81L4exhtWyph4/o4FD7DTU4kl8qHU3ktAHrrzYZ5t3MdwFuqFMfTsXEr4XOZ2EzWARr0SQfsGdMCC2iGZrbgjettr168ip2EkOfGVy
ydLOtZFbHy/VoR3MQVE4MT30yhKDfB0OFHuHuM03LN4H7M7QpklxfsGW5/COb93c9363adBLQUJdGShLzq/loM5Otf+/egzEEp4ZK+hrp7lIN2Uz6Pxg2+hgtk5u141s
EE23HcHLdahVfRP66Qu1xEMn4a1ND3kc8qM+XcZ1v/1Jwo8VUtm8o1UF4DNXMHpiSZad7sn0nYSUBsVZ0IpeyMC9iQ2hLjf/p9Sgqc5GlDzdp6rslDCwv5EVn9IS3CPR
AHJgYnetRbFIpFaSqRNcGjDNOswLA9rSdRp+HZAEsDZUnn8zoLI4AWPiZAbc0LwGuKq0GQ3MFrow3LsEfhVKFcYve0jvJq3tL+g8PcFB4ETsyxfF+E68bALB3tvuoVWS
rNxXNnO449jlyIg8QTDjH5hy9p1Vv7b8HCK4cxENlivhxaUNFttk2aIBExzEZirRN4GANihcbAXJ0dKQWXqsf8UeIJPyHJqcHpTZB96/AJd3+tbArpXWSXJKcf/RgNZH
uQixL8Wig02/+q39+cfxiYFeuo5WBozyp5Z0FqsmUj8B13kdxgu44M9U0jvoW6xrHHHF6GUhj3OeYsOkCUBLUVwZubBVuaLM7e5T43Wsl07zLJup3x/2Z+xjdyymrXEE
+Gjjuq7vgWkrU4KBDwjyPtxImX/BXC2mWjlqX/VW8xzfJYiwXLK2R8jgIt/xWyqNJOnem7AJEo/2i6l41aA/DBYNLb8E/cKoVuh3gab8A4pC/A6lZpxzG7z0vxk2DTPv
POu8QeemDNNBELFb2fPQyMysPdWXIXfbnMTuZkxcRx3dCyVqi+3kFjR+oAMRnMvbmg82q5CXRF3/SuQURTiCPppDgxWs+SPaWsDOXm3buL3eSacSAeHjKjLvlVdqIOTp
b+0or+mQNWvIc0/jnFqsT1++LbU0PCDwLKswDQojSY36TLFLJ+yyQO74BPkD8/Pf2sbLtwZQVACjdw4O+N3W2Ti2EdCQTMv+bep6ip/KzTlW+La36arYbSH2g6UYKCFd
5DETDKdnEzhXsEW7W/plQ7YUthFcjMcZn9ZYGfrXPfGh6Q8tFe+Ok8ksatPA2zQzXCVjPSqsxKSdN/0c8PhDd+UQSEykHp3v/MspPBJf8QDpsJ7uvHZ9QUU3bLsbAIbM
mIgGrIf1ao7+lFjUweNHw44LzwAFl/1TNGWdpRt0dRcb3Ujb3m60By91q65nNTDBgDo+WUbukLr4qlalYUlZLGX9VBo0m6L4lJyY1nfJO6qCXda898m1YhEDDV5hJ5lq
sEqGr5FwNzh2VRv7OHmwmyFztow9/X2cUqoag/TC6ja1KuafV4FmfYbXjV5KfLfDp+xti9foAZfBZ+TcFvDI2jEp/j1JurBDnuI5wkyNleBIN2Uz6Pxg2+hgtk5u141s
lm9Ryelgw6weRxbWaJkYZjwi8QvUB54wroc/3VMIIVcIY/ayIZ2rNZWaw9pM5V2nCl3Kx+njVI9Z6Q63myevZ1K3BJgpWT/bhvqrFVsWdpvDL/7iWLxB+o/glmVt2c7F
r83APINGrw4+FKUmd0QO3uAtjm9fBTXu7oDyIowsBTpe3PZ8VpzFQsHkV6MewP4hcnDxWPaILTh8fM/7FSib6X4w448kgEEoL+hMvqSo+T+zlbRPVcDo7Pcag1i6Dgb7
ySuhJHNouUP9a2gybmioJw/TjfmCwLyiBvkdI4ssWnOKu+t8sbYADGua3ezHvns9eKFrkbXu3a2kjSYfyVivHndSajrbN3jAXSh10H5MZ6pr03PWdkO007tHX7mhMB2N
Cjl93NgwFjlzKG4OKFYQK6CHQqhQ6rgUr1//+zpO6EaYXqbJNuvD6Cl7aZC3shWidg7rETUffUvLyi8YWtUK0g4iyGp46YBC9WquLxBirrCKFpgY1farCB1i2h1/cHri
hVL6OQNCdi7Qv8f3yva+GUUjMbE7fjgGzZVuei8h52ZwO1hbbWDVREueQDInwxTZ8XnGUQJ+Ja34BT6ldAqSc7lBNZJ4F7BwWrzmgHio1HWGw4kdj39gTWoZ3sVyYGu+
pw+DgUk30lRFYZxGhRGSx8v4/2dNbdhbegn/Tk1+LSYNjYX9/w0/Ur6Xhg7QFJVGe8Ay1nLGOMXoVesP61Vq77X7AWThkWAEK3Yy8h86G6wlOkw8blqR57XUoT/z3MZI
DhFAN/EDuncpy5mqY0OHCbMgUIUpb3uqSbIvycL63TEGF8Jq1gO4ThxBVNMuvNaiBqNtSSmMDBJiwKY0/NaMCsM4BQ+JACkMlSumf1qefZTqC03RG5mCs2CT80qz1gd4
gGJxSJPsNQ6L02FA5Irnfu9gttVqOqQM4Ttv2RhoQxUZivGNh8JrNLkYTJgmlLOmmtJu2HX5tPEIsboy000TNnUNhDWCf+SWpaVoV0pQCRDrPINvB8M8Q6HDo+2eh1Ni
KN6XuvdjGHjKiWju0Czq1sSE2vluXKrXg3Hs8FK9SSTf9fuiou42ojzkT4BoGeYz0VZ7777cjxqkpZyKQUj/rI0Z95+F/HRloc5yvzYib3rW+yPjVjESl3cL3lJVFEZZ
JJkPyJxyLJT5Kp5mqL+ri8y13KeJwLIbOoWXS6NmoT0X6Ml7+BZS4N7c41qTW+jSFRe1djX0pHM7Z4j4Xv6FvoEK1IKUwQWISTbZm0QIzkd0m4EEG9mVJ17dWE5OAOZ/
XtSqeKns3+WiPruIRt2RLAzIO1QM6FmRaXMrVEPzPxBgzX11i9KEV2HXd74KYDs5WVs9wj19QgvuxVni/+nCNBmChxXUtBrkIWJC1BLzYMej6BQb8eFVv6S8QgmXfjb1
Vmofedh8EgdrKRNYdDPYcFCZE/smfOJpGqWi7a9+/zPmuI0urS9GLjlMtyG6xFnHNkLDm+wPeYCkBmpG9y5iBh0PO8KM1PvuLY2mOQA86bxAOycLx40EyzLtRpAk+ct8
0HNQNbrADMVsZEyHD4jzBu02jVOSuRPpszpohIVb/iibloWue8Dcou6t7+azzWkxZI2+6MJGwutF71SRzls8lA/BCKpG1a8AdgSj/qW2VvTARxpHQqQRFRXPmPVdte08
YSw6kJgp8rjV9QAMeUWJppL3VQbEhQTn5YLb03BgOGXEmBPSk0KCZ5KTVBLjAZeB7jyTGYS0NxCh537WKrGLySTHgWgbofIaCJFJmCNZflFvZz8WHCAWbvpxrKsuEkA/
wLMVkdamKbcuokNUTs+DQz+kWvYy5cJVDa0+OnSfFn10DrulIThqLP2yffINauAfWWN8RBg5PSHolBbZ75fwxUt7lBmmTiDxDCpuMkb9YvXk4jY5LkIi/P9GBzSsxQ1w
/Yk0QzknxWMZxb3uZsO8U2SNvujCRsLrRe9Ukc5bPJQiQ/OI1nh49AH9U+sq5ZtkdJuBBBvZlSde3VhOTgDmf+QD1v/MjEPXlxb2KM2EzAKTMWYQ64s4weXVnVdlYUv5
bTJMXReM+ZyqIqVoDu6X/4Nb17ftezYOZdfaW9clQUNrjkBAT4K9Fu0Qt/XM+emi+jiZPYg9NQtMVcbpMz8VCGweN5wKoqCU+AM1D64iyyqn4yWFhTgD9fMgdRAuuvOl
he9Ec983yo3jMd9gKBogjPiv3NF3acHH/LkSjCNAhmS4ma7KzXWSB0mN/tJWJOKZEtIqpLI4v3xnlScBAWl774Fa5n0gGlwETtWVG/jMGCMYEzpX5qXbcwqNok4dCGbQ
MfmS/E75+i8eYgPkTrhFziFFYExpEstrpWn4tLw1hZMqhH3zI9p7ws5QlkvPPtUZaTYBztem0/YbrNkYRTzQdj5cCT1qfnqgH4JTVkbsj8lEdBvdSXYEU+mpX0Q8OtrT
zRqFSenvVk0sY5jJJpVNhO4E1c2nzmCsFvWf5+BptHgqkVG98WQv/ozHexdktIC8Fz8JP9zLH7VCJUW8SuPwCthOL8QWdCpgKxcK7XxuHi77s96wfYaO8JhZJPQgsAcW
Upmf2FM9bes04jD5tPGPmpJ1XxYpJ4CBzJILILhMHsexOBLlY0oTnS2PM1HjYcdlJjnnZiI0bF9CUwbZfyvpB33nceTimtr3HBxD4RKP9TCShFEPum5NWjpCgqaDqsAB
+X6rldVQzRucUglMYC2rNgvl4CRvee3fbfkiEGEky8LE0AMscUyBA6tyq6FbdyNpT0hr39G6C7Nbl72rjFiM4k8x9YNsL0of5ey8HHN6TqgLLaCvDmbZLgWeMkrVV6tM
PVCDyX4xsZtm+KZq2GF/iDkOK4BJ/cKdJBgNcaBvX/1PI3V3eKT96Bd9DqfKEWFTogskAPNmdtzvrbjNm3JUyGRC26cd2u4GJQY/7sIJlO7+MW3SpLkoRpOuGKhpILPN
Hy8zYpw4XH/2iv7K7Zc/rYUGIbsTSacoHhi1VmJTDJqiCyQA82Z23O+tuM2bclTImHvK2wxG+1/Y9XAkiXptXZDdT2rcUC5+gEQ/BhhH+/XbdmluBXE1/HmOmqIVEUJH
KkHTYLZ3eFVgR6Fcq8b8rIa7PqTYgvHv98FUJ8Said7e2DfolkiNM3wPtVD1H9Wy2j3pAtgYpKfwypUScekngR5nBMwLT+sElcLlAqzq83BflvW+OvCAwRxE9O+NATp8
xYLZsdkh+tblTmKThx99ScJ4aVU78MKCa/37RhMQ4hM/dNOnpvU0D4ihzlja69YokoRRD7puTVo6QoKmg6rAATj3hVe5QyHxf3f8DitdDxNBOJ8LI7yMYj9UDnxl9pJQ
Fi518gresdGI5NiDeb1phoSikdO5DaEgcbKNS/yJ+L11QK9jDECiKe2yCOypR9DlkQbEJeiz8a5Su6JLfydyX0vhbY7RSZF4Nz1WQY5kQpUJd6BZQdB/neBwyTQVSNEx
U9g2DzTiJIILEZT+sGve24EYwSnT37zzkepX2/YFVBoaRzyUfRUvhS/UYVCId9u3C1gAHqeNtUNUM1N9h8OIwFLK4TporjF/5biAL+PYjZyLtGD9syEqssNvAVeIZSZs
8Ex+QJSeWuNWaaK1wG812K2WPl3UpB+JWOqJkkljU1c+jLMCkituMts2u+u0Yf9yyogm0Sa9h4GMq195YwJtiDiWdlTEm9eTSkEM+G1njtseZwTMC0/rBJXC5QKs6vNw
cQajGhChuFI4IIK5QUXBzbrEjTftB2yvrbblOL+4ekutlj5d1KQfiVjqiZJJY1NXKsE6J7yHb0q/N+Ch4yIKxsqIJtEmvYeBjKtfeWMCbYi+odcxd7veSuvvglcSH5dm
XmPX4eftzVVIjwH0ttwbG3Y8j+sVJC5WMaCFgUJOE7AC6FGgqx8aVMD0PwwSxtlVZ6YqO7UOX2cbWnLGVDUR2lMlbY/xyuTWnMtM6CfKrKLQNLpDtan9hMK4WKfoywsd
LE3lJOD8Jgn7o8hMyX/VhDztqD6mg10pn2h91fPw+xzyPgv7u0TGfLvHPoB1zv50N2quGejbZY9MYqOSJE3RUDDZcYHB5nS9lkukn8Hk2v8GyVlVQDRwi5IfGQU72lEs
3DXp9Sv/j4ac47C8pJ/C82yfkq/wEajxp/f9Z/ZqS8iDF6wa+WsWMmECyhDMlGmFvDP5flkcfWpqOcf0gfqEfVZPweU4WN1j787KT0r1OF/UFmQAXEHAsbtYKX4RrucK
Xhs4xf+7ryzvpJpfUkZcW3MdgO6ReFtkFrF+vSkeb138gCwHOfa5Xe5828ppB3Su4RPLUF2tHqg6wR9bhtCDcSFDP+R50L3e4LpaqPPcs2RwO1hbbWDVREueQDInwxTZ
8Ku+BqLjnoPGzVAlVCNy+N9GDV9kYsn9iPnmYCoomJGcO9WdjnsusKvWmgJT6vI1pF7BopkvyV1NJwXhAxDmPjyJjUVDvJRY8vsblcv0ljsHyVFkGh4GxZmJM7psuNwy
zRVcD9B+wy4Hu5x4D9voaBapRrtzbE1vQVK95IjrJHcaVQ+BfHSIpL0ycoh2CjMU58zfw7mPnV9/wj8mC3DXTUaZQ+JRL5SRviIQ1/dPAAEyIDefKfW5q1v5/Uc6AmsZ
U9XzHZ8xTgpnAmcBM8Y+lKUKo5BvtpFYs+lmoUofH6fys5fFhpbVCD62VXNbQ9Duyogm0Sa9h4GMq195YwJtiLS43aPEijHKvevn0oKOw8LKiCbRJr2HgYyrX3ljAm2I
9eAhsbYpcvuVPp86ImPIqtnghK7al3Gq6hdhkIBdF5vKiCbRJr2HgYyrX3ljAm2Ile0M9wf5cNi7XCslZ10qczoRJszUcoSUPCSCZ0rFc37TIZGc9kTWzrYMDyDvnYgc
P2zHQfiwJ+Q2/seaHkeycbc+P8EqRo3qafd5QWWMNpREouaY/yyNxXZE4AZBmEYk3mmgTjsMR9P6E3+H61FZHRqE7k5JcIxBi8FGWWlmyeNmJJqmAIUP4a7qcx4r1VL6
BoMiHPw5GySYp51IAbs4wWa3CxisC4tR5qTW8kjSgrLKiCbRJr2HgYyrX3ljAm2Ig3EXTn58wwiGNPL7MS7te7IIdzqyNnLRqjHrTDorZj29qJo1YGUl4ZsPVuT9zS3L
z+ObKmeGGpSkXZ1lDJ26mvhEBvR8jhwDlz3z3FT9G3Nk/LHF8zgMsD60bxoHmR5XDgiJKZRqbyAGTCTJqnD+C5KcATrtuwPhUoiksiCNnhawAHQEw2KuVTmV0Fv1Pqs+
lySDAjBAh02hrdKpcENlOB/YmI6aqAPPvs+VhaekZpHKiCbRJr2HgYyrX3ljAm2IOmcBZVUeK8oNMHDzLDhywS5OyyI5f3d7WCESBMS+v1X21HppOtk/LfPQW1clJtqC
bN3LYV0iDCpPt9OZDdfkb8qIJtEmvYeBjKtfeWMCbYg6ZwFlVR4ryg0wcPMsOHLBaS+SnCXsc689kTSD9ABaE/bUemk62T8t89BbVyUm2oK78Tk7k22zoWZ46hooHGn2
w45CQ0p5HQ2Rh+pK9qk/t2gJ3hEJQOKedgnJIfU2bkvkHAnmvR2E1boXqj+Ct1lpOChwhrvOT1+LtITHLffs5YiTzaeBQzdz2bF8pd5cNDLTIZGc9kTWzrYMDyDvnYgc
sS4gW/CIJ92oGoaDREvBRaFS1Use6gdfzwjmLWQPeU/J8PgCLzYC/VqdgpdS9WsvshPhJeOCrw03Aj0EKt7hDqlRFYilDzJ7TInlYsiVdR5273WiI4FlLzoxSTEQscN5
SketYQ33hp297ElwElpQI90LebarZu4zq/2KVy0IDfo/+D5MMUYa/gBYJKGaK+MFAcs2jVC8wcWHV56OheD1S+YNjl87draNXqdTnAgS4LGCUkWJVBuOdFuBXoVkXMox
IDs4j3RIMR3ZgQ4KhtAiibl0PSnHcccydPmXNz0bgc1tu5iyAPWLaxBN9NsBJvF1A/W+ogXZj0rgH7UZrqCCYvvbrEuO2Uwo49Myzp855ykrxIsSAUpSuXimInHrzKo/
ZLoKULp7VyCcWsMA1qSvDzMlm6MZvUmOhSHJUQqQ5XyKDunv5kxEeELO+mT15JIu/WvoYStdFF22vF+PUXop8kH19zmjMLt+en69PwZo/cK1bEh0tZlKOO2AUzAYF51V
0Z2xG8tJx3rAu3XcGVDHalZbb9pJxIZhfteloYiE3pBQYC8xFrfpLcjo2fKbxb/0vy+ugpulqBx61Y1iiwkM2DA04kbPvbTrpSQQgLYPmGNSH07qFaRjO04IjAIz1EIV
O5evuOd6RmnUTAskztiB9EH19zmjMLt+en69PwZo/cKBS+/AVYP5bNK7Kn1LVm/Y4E2qrO6kIiaOWJukSYLg+ACdOaNWWhjT13QwyMixRZnFlrvJj5NGKo1QFowaSKCv
ayWnm2Ga/is5ewh2tIRAW9ucHxc3HXaKmsjHrvitPIp/1lVOw0b08sMBygyM8hNPkYFvxvAeEyhPN/XNmVIbwLjwLm+YIFkkGfi3b9Wyaqdl3NLqeFjXfofRVxzykKou
tkSZP0UcdnKnNNuxKhXdkCeb8j59MtV+5/YovBktizOJ3F+LXX7LW4C4SEkoQKcV4wvC5PjaMfQ/Q3k8KV414KqFpJ4M0ABMjnGDo18U69N4x+kSN9f0Hyogg6QMSEp5
xDfUMBfOBQGLHobut5ZOPhXslHzqGHFz8k61VazVHKaI1k7lV+t7PsfkeR3kDMEz21MGHvwDcboGPUZOwMklMmIPbCeTV1xGzA66WlP7Jrvtsxi/S8JoyAA4rNLtaLak
GLnrUxCwy+g1Y7VUr8uHTKrXZUUn0BCSqsD4jGydnWoDW3YYKRh6K6k9ms634LFGpC8ysLWQq23Hqulyer6/HSNVGYetirAz0iankvDHzYX44RaYvq7rYwxiPoxnwBUV
9iUzka6E6+g7s5lkZ9i6hw4IiSmUam8gBkwkyapw/gtIfJLwI30qbKjuXz685Hs/C2RrAtyzX5Is1Zk1ZcX27xH8X1KJwUC/yxbGEK2PSXPRlnDCDpUCG+DyNddFXEcX
Jr/rswX11Sdu49Hu3Ueb0o+nPegr4Cxl3jXZgN1AFZGAhND2kOrUdfrhQQUK26ywa/V0NoG8Zly+LJM/1DDxBoEz6k5ZOdBxK/ELzwLUeo6y10FEoPZyvLxRLMeJE7nx
tr/t0Fn8rzYf2dlnBHDVJ4knfxXE3zNJAn6AFbBQgAG7sYxVhRZPMo+9M5nUGxTQV7h4ILOiSORxNV/TwDa1ZnT4RUb1sfzm1lFnsQ2JYsefbkzIUEJ8x4LSbNao6iu/
+YEgYFEMMlJZz5oj96M/6ImP6hIoQaccpBOA+3SVG0ZVuRCSSo1/GOMrbnKG1fV0AkYMjM5w4Y569mgg42Z+B/faxi4zU8vP1KioV7vD+acky66KRSHkipxIIVJ11QaW
2On+Zy5Y3kYCwiZ/MqIoV5kVzU5nqBEyoyaT47sLoQ0xXlmdtUZHH8CwB6dtBACxnzdbg1W13yhLRHUDPEEGr5INwQ5HcLBzxbbyIC7NgmJqP10fphijSeZXZORr2Vwk
4mQ4ujGE/4OEM+Us7v0ao6QhMp8ffJvlqm3PsgRVSMpa2PsnsXs85l8sB+pnifwTr9Gfe/T8JiNhRB1T+3rGSMs/OmHXakbmwxmhQAR2XNyoHyjLQDtKyHhKA71uUJOB
B/sbDwGj58drdrTbRRvt+ySNADV+7I57ZqFm1Jd/fQ9tkXPteJZX2bXvtNLt28qhmudFA1A1Bq9U5pma7ziM9BmL3S3iXxS0kLxlvC6Nlb0jJohzPWpCUlDRSvWQWpE8
/Jr8P3eeTB8JyzD42l6dh0zdb8eCngI0iF4V29iUOIPgfFUxwaBf4eypiY5qv9TIohakS2fdUebEc5dXXzqJdGpHW4VoxVWGs7DLrI9FNAbr4FaDKGK3FhX/0d1J9BM2
8dV0wtpfk67rR2XgvGpc6Jay5x3S4WsuUrUEZA32z20ELcp2URYmt3m8u01wVX/jkecl+LySf6shJkgeSI+Qozift7V5yU0/1fJ8Ra6r3xCIAVMlZij1Evtq7wYIUjID
8J+IofKRMEdC2Nq/5EJQX7t1Gbm3vvYd8asI0R2wwOCcPXlZT/zlkcwGlPP2z0ugnPWTWmEnOkisY8QmE4r9vo/UjJRbdwcT8CnIP85ihE933CrXtnUMpcfOzHzhzpec
xpo5JBCNPQ3+KZZpFFh9dFS4shrNqTAu5vs8oAaY/dpAdVYtKUdoFF0hC6vtYuEpIVbaraVCQN/oV1xANZIidspwAXLn8HA74yuI6RQairid0U2fzFqdXddD+9SvqPWG
ZTAz+NYkzprrrxAr2c9SQZ+BrfPvF+1dkWEiEN3tiGfxUEsXz8GyUTJuzajC9ZqX67eQYgExxubZHHjubgvSKY9Z9Vgl221/xo8seQ7DPJi2hGXb2sVLDhJSGhB3VPg6
961Kjjok0iHYUyDIOR1YrhIY79IP23h5mKsm/QBLusTF1BiUHYMS3PxvNiqYmh/HNVrXyY+hOluQlSqdcQzUPog0gaCIqS7d6ObnQzRmu1adq5OIZpF/DbM/Q9E79Y43
lp0ya//T30to7GiCAGfd1Y+dQ+MRJTY2Fo478hgxqyCddS7m0N6MIUjcWdyOeVvpWW7IW3OSnBdi0M51cdmF93YZ2dxyLgnHE/WU8Zng+U13XDw+5SeqU390FqCTk4Gb
CPbinw9DPq35tJKxxeMhXODVFITm9YAzlJIWOCoHWqTfix/GTSR/RoEXGo2szgUTpAUejK26rInmFr4gzopwixS50hOXcKH1dB7Tw1S0TJWlM5A47FhtQ0b4YQfUsmEb
kikicTixje+niKPzA8hK3LUpg8McpF0JM9m1u7qpDsXEBGeCI/dIgBD6QhNCBSLikakwqHi+SyI0Tm8iLAwQ4F1/Fmtsa6zuUQcJj1zU6MhTAK76n3Y9TjNbuDrsC6b6
d3LaPDo+X8GLcMAazmg/ACmZ/Rq+xq8GCneM/Myzi7ThFXmAbR6Le3mBWzt5QYgBd1w8PuUnqlN/dBagk5OBm+2jNpXFmceod4ZEUzNlbXla6c0dPlTtn02qWCQADC75
G/g/l5g1iyaDAlt5dy7BoPHBDd3Ho/srPa8c6tDR3K8m0EAfrkUhjoKOvp2oCLXlWorFZiZ2n3xSQOOaTQ1IECj6uxnIM9PTrWiAduI+c35HwDTaE+MBSftK5YnTAqIk
a45AQE+CvRbtELf1zPnpoj5SUsdmjor6yYIb6/mMt1LK77RB6IEtqVOQ2ENBHstx15fuaxcRH5glNRMHkqkZMg+Y8DeMBrcsdvweBHO9VuA37ov6RDpywu9Vbqv+ig3a
Zb+oC1xd6BHN7vi7Q1eiKrBn0DsEqNvyb6c5z2bmzip22bB/OEKFyFKHpSWlV0EO3pjliHrpPXHESNW54whttZGUcu2DwKEKLBjC/Ch0l+UuYpGIjaUi7tf3s84xauPr
a9Nz1nZDtNO7R1+5oTAdjQ+R9iWCAo8oTGi1r8eMhzNgzX11i9KEV2HXd74KYDs5S3EWLxHzXYETPjwjPxUNcdkUkRhUpu1xxYYmXZZgJO3fcc7Uowv5v1vZBzf7hEc3
EIks5L4eRsP696OBQBRhwXhUw5uTkKx8pCSA6aHI91IecOYfeFy8lI2Uj+LFvOrIy97AUiHM/DkdT02yVCIvljdm24RxZXn22iM+8LCY0LrvpBLTVdQHkf51LtYYmUEm
32dn6QvycyTFS8gFC08DoLh5w6FPWC8ZWQNoWB8q+zTbB+w4CgwMmJl+OIJsV5/z7TaNU5K5E+mzOmiEhVv+KH8VWtXhybXXnBg54trEYvsk8Ks9+UX76NA03Bw7NDhC
5OI2OS5CIvz/Rgc0rMUNcIN7shlmSZMiOFEZjYooGPb9gGLjbMRKGA7wgaYnUFPHT/19hnOrOpIsBKGhV5ccjzSfjM++WWV2URRVjJBZb/dShpIHg/AIpZ7VhUJ7hkw3
Hg4QP4kfMxTDLoOroOukgTs+FcowHIPWZY/nMBcBQ16QSAAnh27ZyCh2gK+b81DdWAX0aSq8jdPnfYofg3WoHRVC632IYayIYTEgxKTAJKkucK6IgPfEkwHqN2QMFuDI
5XfN42XVmXs04BAlOB50AUAyFOnSfcqe6PPzdyRxrhRKYC+NoSJyC1S+nXgiLYpJDxKkiZSl0Vk6HLEi3RZhrNhOL8QWdCpgKxcK7XxuHi4A0jsNpYFL8tawNXiJJX01
adoILGXn/Fl/Q/i1lZqn180ahUnp71ZNLGOYySaVTYSPygrp/RJOwDAsDl8AaV/BK8SLEgFKUrl4piJx68yqPw/zsJR2B4pmizngNbXn7iAQYbAbCwlSpiO7mxmF8IjY
FpG84WsQo2M2lW8CL7HdIRrleSWU4wHkDqeLnCCLXVdHbE8R0jHvFGkRAPbPyPGBxOtZEetHIdx23QNhkq6QYlkJrQ00tLgrNHqy59lHZ1BVnQMFfL4QuR80yQcwzKXj
wf2lfLI9xBML1+Y6GKcQuRE4roXEfdPzmg1vJfRNDNu5/wpvuZxdMN+D4aP/jS+Za1WcsKHYaDTx+M+18fuablSVaaev2TpNch9HfYDz/avBrwZZAbTiws17NmKj98u+
pmb2iKHJf3WzPxNWzCtDXwqp0pXlNJI1V2Jz9InprAipBDvDR+r6EX7rgG6WCjXHCxOq8gH2CAIjlgGbrcfcM+IePStPGhnptG5vwBOv6+bfTGQmVTAc1WWBgJa/S+Bh
BJNYoaZYcakgXoS3+/2B6hU+q09ZFqNuyLIhM20Jv3FKYC+NoSJyC1S+nXgiLYpJcI9jJwoDilrpW7/5GUrNzj1JS9xQs1VSbN4vF21Hb41939AvFB2MUDj3KpsFUARm
JsAxv3QMdUIezS614N7SaKXOGXM3aSeieByFQgwecxAv/6ECQPd3JzWY2gHZDyXGkQbEJeiz8a5Su6JLfydyX7QMf+xXJNh0r69qpCM7xNGyqkQLdU7I7Ms/gP5TrGUa
pc4ZczdpJ6J4HIVCDB5zEKOVVJFxi6uJFJLmX4ahE3quyCcH3NKNi54OjWYgXTg5mzf/8Xs+u2M898QoitOsJ8qIJtEmvYeBjKtfeWMCbYiU0B4T78DWssZac+BwRkZK
A6EvQWzZXRgKAFppQ7PQTipB02C2d3hVYEehXKvG/Kzsu+XRgGdYrulj7mbX0+Y/3tg36JZIjTN8D7VQ9R/VsovzsVukaGa6N1yH+UEpqbUeZwTMC0/rBJXC5QKs6vNw
ZVtNWlDjWITAoKtmOqXCfOzyZS6xLALPvfy3rhLiu3ce/NdIzTm1IkwhXCricFAzwB8h3XzP1Gut6JrYQ8jDVMTQAyxxTIEDq3KroVt3I2n3pdO0T3dOjuYNJsZq5n+A
N7aHq3JCSuV+PJCN5JOOgoSikdO5DaEgcbKNS/yJ+L0eTfSldNZJReceJ0GQB3qFkQbEJeiz8a5Su6JLfydyX8p8MzZymID8RZcLzQN5g4IPJMVkT6SgGrUlUbEYwLM/
cD+osMRFs4t7cd2segRuD74lSzGkH5UmXAxXEoidWwoVHe+GUR3mJWIXnCtmfDERqjGIckLBSyUcI+QOwD5Vr+lrmS66CxwFqp5nlDzHsgLj2KSvYoMebAYY6iiN7r3P
Sbsuy4VmTxDqVGTUUZ+rgbDBTeDxEofzZY0kSGtPrRQqQdNgtnd4VWBHoVyrxvysqXbkzTId404Akvm/47VskMJ4aVU78MKCa/37RhMQ4hPNCEcLv+oaRO+sdyhFN3+l
49ikr2KDHmwGGOooje69z1xBjiGkpaVxvIQfMxfXGsaHMkr59FzwBRrLpdJB83X1RixQyymgRePt+nY/nn6LzMPP40lll6O/TlCZbUSoBvdLvOI51rvaydR3Jg3OxcFz
DSwBM64jNI8imM3H9BtmU39p+G46I/AjpEfkYZ584fSFrNQzKFxenwr/0FPbbZIXhw6QUNhifXaS5isT2i7JkDJrObhynd/wcsAbE+ysmimO3uJWX0qVf6QyuKQxTNO8
vsXun5IhB+85/c1z0W7fWK1viWE3G/X2tNFbHzWyr+AiplVY01fVC1iV2ck0MccijQ76i4WIddiFsgFZjKs3CrWgbc/Y2chFt8X/Oukl8SEyoZZleVUIaYpVhRldguEb
UIJbJm4r0scd3jBJ0GencyqMxaEmfozb2kfBlWesQUibllUvymDcdXpda2sN+5PHa9Nz1nZDtNO7R1+5oTAdjWYB4gKXLUYhZMtDtzlGLjaqNsyrvLtNNVNBYdXRpkc2
ziHm0Il5ydSihLyDRMER3iIHTB/lhWIExAPxQR2aMt2OLoYGmsr9jjhp4UCidXIru2BL/rRv6BoVRaAF8ZwltdZ2PS8H36DETzePr5Q/YLkFoQKVvhZ9krM4qR8IyaGu
EjxGMxFblT79271EGwQ8BfNV6K2mDuJSroFI1QSq+eXx+BMC2ItF6fUWRXz6dAj1MV3FIgDfvJ7sdHCaOhuXqYplx8KUWpOknMBrGaeLhLsWmTDHZnCMd7pnCvC9IPQ2
ZDKU36+g4qPC8vT1SWHMp/970MMqfDIrerwDWztThaZkpd7UQv+/lKUMzaKaUevleHX+P2/6U/ZrLoRWTC1MXsAVb1B52I+P2UXOcAb/XRVZMEY0bJxpDeiQ4sTIKuAh
xpLsZ8ZfPXe2l7VCyT4kpwAGbzMUslcQQwEZf2DIqlBS05M7s90EhofheSI9h88ag5fbvipBqCi4uf6cvzdikMqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13L
WAM7qMSqR7P4pQb+ZPpd5Ju65phSm8LFZ4YStSKkgaguC42N55AJm93gTOgPDFY5yogm0Sa9h4GMq195YwJtiCmwFpr7r3fIpVdYnA1fXcvt5GZtmeaEtQyyzRceW05Q
m7rmmFKbwsVnhhK1IqSBqKJMY9OHMvThkzLucr2H9BJ/t4SHRrYqTSIrk9prikLIE2G4P3w8HQR15weMlpCYY4tEgQ8e07tm88ELew8CHs4BJOmnDqjiIy9OxAxuSiip
d5Xvuzl4den6Rn/gvVwk1cqIJtEmvYeBjKtfeWMCbYiR8vGvreuT4JPWGKtJ+JatQJEUjf7QB+1rzxbXWUr97PiXj/adrWMOPVpVQNqtTCTRuze7KE8ld9XhJWCImbjI
kYFoYFWrLJNKFol3u47tQfHwt6ZY7te41bjeK9e2TnPfAffdedpGKq1rXSGXjvLas9onqZcWsUjN8gH4tbeOfmZPUIaY8nnHEEtsz52et5cJisM/QUoZbYrqrxnJNbJN
bj3Ko4+CjH8yg9uuGxmZnU9AHUqNPiKMXd6TmqYHnDGQCER9dmVVn/fLq6032MyJAPnhKkMwlqfLjKsd1zmACvbUemk62T8t89BbVyUm2oJs3cthXSIMKk+305kN1+Rv
yogm0Sa9h4GMq195YwJtiDpnAWVVHivKDTBw8yw4csFpL5KcJexzrz2RNIP0AFoTZTZ7Dojf1+m6i7iMb9AEQRaRvOFrEKNjNpVvAi+x3SHLKKgD88PC2+FONBAxWS1Z
Seor+1VsbbG5l68CKHhk0j71HTn14m81fQy/PIbQNkR6ijmp7TPsHk8rdG838NL6TazntDzpZp7xB8xtw7gHPt4ER6ENG7m0FDD1bgBFTDrNXtLtfDARzwmVP2fLjDqL
zryH3oMad/wXhUl6fYM5FICjv0vYGEGhB3hfzRYrxHU4PsN2kBr0hFOZn69EBTTQqAiFsBwMgBtoaRm3YtERU9NvTiucfU/uZhaKRK39Ep4NvY0lxum7Uk8eIn64Y0Nh
heKHhisE2LN1sNwUMKb1YKii8382Y7mfd6YoLhy/KpnR9vf7rICwMQjq5hsCq3Idq+zfDw1vEPfHBe/waN5K73qM+6xFm/p9xJebZoWdwM/UZr00StuqDtIK1nhGPKbQ
7QG9rxmiZY9fytCMX9apMNETuRGb+qODVlTw6M9r0nGCrzMI2HiEl4XdPWMpZz0Bf9iUn8v5WmWyHeErKoRoYE4HBryYQ+SEKOIZPV0CmUlwzivfMNObyYI67Jj1ij80
/1frVYXXMjlXM0POX6fj7dGdsRvLScd6wLt13BlQx2p0au+WBrZ4u20tJKLAOWcQAJ05o1ZaGNPXdDDIyLFFmaYnA/4b0tR+CLSD5PDl1rLPpmEwXJpWpBvqOV5p1SSt
c0fuAIm4KTWJjtMq2smFtRNwC7vDXdezWJpG+B70uWcBEZgHbvLtzYJ7c3+lQrJB67O/dbGIrTfKVmwjBy2GoLjoTAR/pMjxy1W8yaWARdBoOQNpNmVRWX3jnjYLdG+D
AJ05o1ZaGNPXdDDIyLFFmRKHGD0mAo5TQ6wOA89TAGiywVwBkHuhGU9mcd5Ed7ZDnHIr94n0WJE9pGYP9devr5mtWzuIAXU9LoD2XDO6ymiZIHLXJz89KkMcDATmVjfv
MSp2BqfzXmm7wJuM7b7lANQ2l1PjhPyQ1SvLuRhXmDauSp3qtq8hGk1nG5Q7LSewj9ap4me4q518xESU0JLbS76AKU045j5kWZvDajlCwLXmtSvKUuUjYx+gwenIzco3
Jux8z3ndnykEcwaQVjwSsAeSjzmNtFBafnE0LWeXVY/koVkCeBj6rcrtYYd26Mf6wuPlOl6hN29DX90GhbrmVeu4xTNE3WnGNbubyWR6h/BgbMQPd+2bBVsIHLn/Z3X+
Faa7RFdo7DbTOqeRHuARjiSXI19mg7wesJeaeR4kWCV101jQ1R9H79hoZ7/NPyo4qYZLG8os4pCplG/VU9olJq6pcuRCpDuIGK/3926DHQXk7hCbtD7wN6Ko0UznLBG4
dkelbi/eD7CZzNekeXTDNkckUUpJmX8dt8H32bICmuEnD02MNP6vfu21C88h+blcPLh55dlY9pKqf+2oUBJdL3/0M4ImSnJM2Im/MPFffnSaEzNfVVANeg90trISwHwT
3kPHDNyvoGT+wG9FmHcjNAC4Q1tRVaGZQZmrwRo6c6ARyWQDtO5Ej3oaawJqGm/rzUIKZJohsJfjQ8SK5hOIT+1zIgJ7L2c+1XW1dJh1/t210jcgq/gthtIlUQGrdaQF
hfOp3YUbq+6JyOgg8mJ8IfWJ8t/ek/hhBivLpUS+vSKuKDbCpBTxEJHWohDZovv90+P46FRc7F1gT/UNfoZFOShaZC+Hf5vPsSGp1R/1/HHhWJ61y5hGMwMuRSUBsFDE
/rNLkp+UPBt2nSClE9SDVf2ttEFN6Yj0m3P/NiCnW/cganG657ym0BOcFVzH4tDuHkqUZdGHJ5zoeK7Q3gVMVukkVidbj2/ubMkIcj3FU/x8rB6E499qYvgKggWsEDrr
99rGLjNTy8/UqKhXu8P5p+2arMM6Z7SdBcVjZ1u/JTI9x8fAaxOROt4e9IkO23uhNR/MzNbjumL21INUdvKPUd6/2kAFYsSLq8Y7tuOhWu0DM82tkuzbcnw8jGhHQRBZ
r5q0X6d5682A4jFms8o5+xCG503OLOBn9wAfhM75DpZNfUbJm5eJegNiGKBp4wNEnOwPSD+ruyNx0Zlc07FpZaHHb+Xemb7SAhT+BsDXQNDyHOSb9wD0dEvro7+oUcNO
lM8QgaEpGtjuLEw5MSeXASVcueSzVmspUL4IKdM5OOsHVQexRelNOZ10ym31b5m4jXHhU4K+IV+NktwNAxqPO8KaQ+LG1z1NXn3rIGpNo9z+0TZDdDlm+39VgPCwBQlF
N8QVsEnzVC81c4W6YNgk7XUVCRRHe9GqNXQ1daUW9j41rjKOGnqdieuQ1uzvHtZMxHfoYinCr9CASde3T47YaZ6SpsHlhEuEhPfSFO9ghczVXJwabjUjpEYXjqFiv85z
P8rQx0J3P9uHsYYHY2Z+1HthlEdWXe4N6twnbXNN209ELjKFmZzyN3/V+c/dROeByYlbupsXY+mzDEt26T/OZtxm7fN+t7BxTFyzPkp7gDtOnSq2dEyDi+8mXtLpvHz5
l13igCKXFtuubJNl5OdJxEkmLswK4r8tNFfSybJsSLqlZdEDJWWDIhHZWRRiDULQg7tiIrG4XZ/cqflC4/3S+rax1NAwQoabQF/hr8thFQOKzykgVFIyB2W4K/bX8l+9
sDeLsZ6K9vnjoyWe7ZgDyakBp044HoXS6ko+um2OtJJyyL4cM0dHXhw+JX+G5k6JimXHwpRak6ScwGsZp4uEu/YXpGZxuZHlEwFfHqi0DjIZ/FYUalCpgL5ethDm00bW
PMVdP3/wwep7+Z6U/kKzznIw8sFq12wWZpq/WRTARN8it1Oiqpt4IU/UMM/XipR+cjDywWrXbBZmmr9ZFMBE33i0J7DDvlmDP+19aRGGdYh7FyQFzf9yZJOT5VgF7ekF
pU9jG2s+QQG6k0tM+Gi0pz6tjTFVq/m8xRW6j8zdZw7DdBdA1kvYY1u6CsSRa5i4VGGAfQbSGr9o2lcpZCbKeSlnsKFE5LCIvvy3yyXvKn85tJcEeZncHumHaaKxwYSN
4dz4eI1Td7XSKiK6BkzfKzRWpGs8SrYPkLkw3kOf7OlTAK76n3Y9TjNbuDrsC6b6VTXFQn9gqqM4ZHFYSIavD0+WH8P58PcjwgtbQYLNVouIETgn+VoGqlluqCcEbbi+
EBUbGSMPtTV795YRIhK6b6Qtlgvq5Hp/YwOX8NE5+nkAcmBid61FsUikVpKpE1wajXME+RMUZidKNgjPXTJrUIzBkSc5QeW06985u5RToqpILLitZymLc6jHKxj6tqQg
PifFznQ+SuBdgStlL2zANZpzasvwqpGM6sFXbDTqDkSKNctimtHsFRTeOUzqVNtJdNvNiCvIDTYZ3TWNOyXDRiFW2q2lQkDf6FdcQDWSInbKcAFy5/BwO+MriOkUGoq4
9eYUCpyIiT6viK9R5oaOzeM8dD/fMH80d/AuBoDPS8NUYYB9BtIav2jaVylkJsp5nK0ASI0wGxufmfA+4jeiq3KNK0IuL3KOQwKrCxaZPQ/j9raXfOWelmEFVaXO71Nj
3o2ueDydH3fNyWgCFHEU0Zm5SZkaklWzEfEhOn1bcQadgh87pR4YqJD4XY+De5Bl6snffk0FzjR6/SlHrsVVn+hdtTRBIr0YN4IFF6600+6oze0/q26D+9IFve4uIFxi
jeRBO85tBVCTXxvz2LmH86Qtlgvq5Hp/YwOX8NE5+nn9sY4AVGrovl6o7YI2dGhiT6uZKQhjnalckN01lGhQXfNz0DVK9dksDoV9OQh4idsNoLFGfnLasQcS/2kzJmqL
HFMVXLkE/BKo80Rkc/Epuim1cBb+5ZiBOPNzcYxHktHtNo1TkrkT6bM6aISFW/4oKdaYSSvzPuitEFuD9PZeL4W+zQVDCQI+Vp5L1FXFLj0kRB2qQSb0/FGMuyvYndUr
og9ou4elbXSr8LzbsIrHbXcr0XC6wFHpGpsvYJDSxPEWuqSDITS2HARTuWMq5gUjbjFWSJsOIS68puVL4ooWgrb1aRqCVh50WBDzhlIeqeVr03PWdkO007tHX7mhMB2N
JKPRxpzQvAliLamBRY28upQnUhr1Z4F9WrsQBhwNV8Br03PWdkO007tHX7mhMB2NQDImooa4QLxzqRJp+nLDltEfIbWK2SSWb4l8FBlJ7VJel3MuFSIraOKu55trqdsF
36pfX4Ld3/KDRRr+7E78ud80ANObdtyTT7AxPSmFQ9+3fMNIUnpqaEKbyfzHn0O2WAX0aSq8jdPnfYofg3WoHaBgP7bfcllV7b5Vg9ybAqBb6XPlPbiCW+NKOZ38kili
yu+0QeiBLalTkNhDQR7LcT1VABLjmbuwDUvFNfIXku2jE7+JbUAV83FXqx6D5973ADzOLRIyu4mLDebjC4CN/K3XZojBJkZuxy5HaO5qEc/ftTvS5k8jzHXWUNfjgypr
Ln2d2Ok9xoyrq4KhlSBP0ha6pIMhNLYcBFO5YyrmBSPCJ7zuUa7vFXvHFusKsHz8a45AQE+CvRbtELf1zPnpot6Y5Yh66T1xxEjVueMIbbWQ75igxPm7goXebDOen6WK
a45AQE+CvRbtELf1zPnpond2VV+Sw2rL1xRsDq4B3mN0m4EEG9mVJ17dWE5OAOZ/1CG30Lcz6hZk09XfiZNov1ObH6yLLgULvr2D9+ptfVB051SRsudDgGXIrvjNUHGh
+UaZi5w/xQrMcnOMAGc9JxCJLOS+HkbD+vejgUAUYcGFULktOHFo2ar+AtXZRvVIOZeRnJhDDIn3NvcdMl8guiJViZ4LhKL1lWTc7Y4MG6/m7HzaiKUDNndk0yYS5QRr
JGmmksZIHfhdHus7i9/NaP9+Iwi/SPt6VedfFOTCa2KXJQeK6yRv+mE40lZZthpm+sN/dqFLw7yUWFQrd1Ehp0jQkG8le/x1eKfI44GXbX4S8CZBuyBqPRj7gKF6Hoa6
79r5D+xSSWBz3sb0ZSk16ajwcPAi4HIMq0XZXN4A9rolQIQUfhNc9A39rHziSDruviRus812Yn7eaN5QLUlfMYlcINQm13n1gCgseuv5Q+cTg67DDWOub5JzztLJo6gs
xJgT0pNCgmeSk1QS4wGXgddXHP5NHhTCaMwz1mEm15EnaQofxshAZ/2Jhsg4GM9+cxryEcozxNSLhS3YDpFWNo9qLs4M+FDeeB3BuUnh+BnGBl0Gd6IFbBQBvD+SboMX
wrhRJevdPwd480hzB5uDQbh5w6FPWC8ZWQNoWB8q+zT90yCY6vpiuHXMMrjlUXTd7TaNU5K5E+mzOmiEhVv+KLRAOKhxgIprtfSzgf4qU95B58nPzQkRw9xA/iA8ZTYp
oVUg6+gcBFVkYyJJXiA6R7qWCWhD+Q2nzNtk3tV3XD6GF1o8grkSH2eIo1qVDdA8eRoPv1ello+w8rbx53cSB4ZsqCCPstanYUe1+MCusrMuYpGIjaUi7tf3s84xauPr
2GtYAYWDc8z7u+8JeeP0HGuOQEBPgr0W7RC39cz56aJ8mvQYr549wFMYZ7sfMsp7m9gTYeeU0JPm/IMCBezRabbYfOn9u/HnGp3rK1Z6NxlH6xOxSuYx0DATadgRE2i2
gBUXChQW4jk9V/40iULYjQKaDQr3ddNNd+rwwi0/p4c9NvhuYFx3mUy1I0bfoLN8IQi7RvVMSV/r+cyuTcIrCAnhRWNzXvjvKs+h0qNiDj0Eob3ZFKeO9kMZQLP2/35O
eP24O2Htj0vBFCHQQGphiTKwnbkZM8pay7kqDDnI4Kc90U79mUrprtn4L6gWPc834M9m4712OSXfksHJdQCD0pwxQyrRpCoKa+cdyTdaPc8CTVH4MGfQE+oExg55IJRJ
nBLVi5jq8cQvmgjH7oWJqaC8Z4OMhK8mwUyzKfTeVrKtlj5d1KQfiVjqiZJJY1NXuxUP35koVOYShuNtXXlK07F70n3BsRHmaaeIB1odgNXxzUCcbfRX9Tk/OflME62z
UpEJcA+JoTc5gSn25PctGM1k/7dBk4s0I1ZMXP+9pJWMn6AAHZ5z97PTbMdx62NXaCM9r0vzWDdoUkjzHnqL6WiK6m7BRICeZqkRFs8bYa+Lkil0UJwP4VVNvOw1v37Z
8qvy+zuP6lPRc8PxE9lQhePnsZpJMc3cfBoBOpI7CZU1ZWeYDlMtzxoLLM66UKf2pRhAsC3Zxpqd8EU2rAqtLVGi8K+QXQ+b0ucrpT9/ntPnyaGN2datPcJmTL20fmGu
Z0ph5iysJKER11Eget6uRcBtYaz7Dj1vu1zbwHr57R49NvhuYFx3mUy1I0bfoLN8Ytqlqch89ruOzqirROP0yHSSlrebY3kSVqILGcEm1Ce+Qtw4e3tAH9xywKhquTGX
R/RDRM+RhJ9jetuFEl039dU1jNLCBwiQoQRlhuekyF+SZqbK2TbpizfhrB0gi0m/p+VeT5e6VTb52hthktH7GEzDoQZLBM/ceqbHDMFZhcttnnJtAJm1sfOl4QlYSufN
1TWM0sIHCJChBGWG56TIXx5N9KV01klF5x4nQZAHeoXKiCbRJr2HgYyrX3ljAm2I/pUYWODK7KdHzx4MJXdLrd7YN+iWSI0zfA+1UPUf1bINNQCM0j8/CiF7K1+BMf02
HmcEzAtP6wSVwuUCrOrzcE0CfvgamVFeeL9aDnfzJYxZiGazVaCZzl/eadaSBOywwnhpVTvwwoJr/ftGExDiE3C3pslwc6YcpYQIOBD07+C+3YqARA3TNg5fUiKKMVUN
0z6yYGJf8gowrWOuNrxKmWdKYeYsrCShEddRIHrerkWN5EE7zm0FUJNfG/PYuYfzdJKWt5tjeRJWogsZwSbUJ+wcp3qAAlEkRS0Dl1a4wf07sSYVHeyYaDC+o9o3Fzvb
AiMcNlGgtOiIJ9gdZpQuIM6g4dPfQVMpC7/Fm+iI15TCeGlVO/DCgmv9+0YTEOITitAHBSNavx6SnQhgl1ax+E728kUeZ7sin9oWLIVFvlNfLrgJIoS04bgbZ9RCK+d5
GnsuvmjImTG225e98AicyNg3V296zJD4Ho/kHecMuU/Tkrk2yHPcXEvTZHl0p4rorZY+XdSkH4lY6omSSWNTVw8RkJk03+ucT0vW4dt8YB7MB+9cadiOnkTQ0lTocvF6
iJ0IlXP0NWP+sd5/4GJq+83bNu0gJLss+nJjcYhLwlcYU+Xz3ZI0ikagqg0uXLH9kmA5kEeVSOFWEptFTqN6HZ7D2Jj0FRffxzCE0eHt+0oNLAEzriM0jyKYzcf0G2ZT
f2n4bjoj8COkR+Rhnnzh9KzHF7th9WQddFai9iWWWSaHDpBQ2GJ9dpLmKxPaLsmQMms5uHKd3/BywBsT7KyaKTd8edO1nSFZggIQIOSwmj/A8xOpUkDeJGJ3KqJEr5dT
u1tRX6mq6anF3WwHjkYIKCKmVVjTV9ULWJXZyTQxxyKNDvqLhYh12IWyAVmMqzcK1Ndwx5OldW8thMrNSr8oR/YGEVzZ/za28jwGo7WItuJxYzhB24xqlPCSqYMisofy
7/vyiBjd5PSTkGU0ZaITqt+P/qMcy7qPvL9LzK4YJcwVL6tN+7ixG75+tdyvXsJrdziP5asq9XUdhbc0FgvbjCfvmQ5wNhUm7Qg7ekEGENJ3bYnkhLwBoHF4TX3rU9zx
a9Nz1nZDtNO7R1+5oTAdjRYLR0F4H3VS81ro7ITY/XO+EGvVB5nS9lbJx8mNAl7Xw9IQsZ+1ZKG6CukAQSPY422/If5a5xHXDcAK9m/3RQ9Ed7Eccs0/OchV8nw4rasL
Qp73BhUplS9xUN2knZvpRyisPM4vWHVeoT+eBLF1ZeLwNr9kQd9vBzw+Vsist5hsbJhJ7g7lXPQmAxTffeqh5rmGYqeiRbYgkdTcz9EALao6+4qH98LHP9mmENFnFHWk
GWXP9mwRR5M/7vs/6FY7qgfJUWQaHgbFmYkzumy43DJLxHEfQ7gaLecsIsZvKe9DEjxGMxFblT79271EGwQ8BfNV6K2mDuJSroFI1QSq+eUCpfC4+pjhXJgPtXYnYUR9
OCFmHc72OnXXUW5iIiI2PYplx8KUWpOknMBrGaeLhLv2F6RmcbmR5RMBXx6otA4yzgY+b8Ry1UBsEUMF7KgmdD+OwPSL5A6aK0NMsUdvtfq1JdO63H9cIw4KZQDJjuVy
tY9ly530I8KxiW4mdG0gTVt83EisbG4jD/FCJ+k9AyiIim86cMuJBOYeVpcZw1W+9c9Sh3x4AEPBLrI695I3QXYc4vkRUI7K/t1mAvm9ulfKiCbRJr2HgYyrX3ljAm2I
0Lm78rr0u4hTqTje89kJLcqIJtEmvYeBjKtfeWMCbYhyBy6pfPxUoXEONUlR82N2awFJ8Z0jw/DBcdKrMh1fZqJ3SiBZNStaEB5FbOxR1/SluGpEylCNG9iJGZ96/Bq7
qWW/CNnulht/rLzYRYgGCt4ER6ENG7m0FDD1bgBFTDp6/wpBha/M4oKZYLlfhFJx7VCFwr+FuRYf6Fe8rBV1iJZ3HePSSCjMeUEJF9LjuPd48hoeZh2cPYhblve2jWO4
vmLIslVOKDuhqvAjlUA8lzkg90UU4jFpnFIN9naT/uxMAJrDHmKVuGFnxqGbA/1pYNLYKxdBjjxtb6GvKOUTFIiTzaeBQzdz2bF8pd5cNDLTIZGc9kTWzrYMDyDvnYgc
OQE6ySf9qWHku1ohe7b0UUf/X0EjSK1z14ghty7bfR3J8PgCLzYC/VqdgpdS9WsvfXwI1US6C8zsPgh8VL6iq6VooKDyOMF9v6ksORVTaswrI9qW7QCu0/oTelnCXD0J
tv45FULL08z224yvIMq6g1hJj/sJC4BD7fzjlccuoW1kFboHxZsy18HK4jR7W0JAsmn9Gfc+3utje65cXRaX6MqIJtEmvYeBjKtfeWMCbYjS9n8LkPi7FXyEZHTrIDFz
qhmo6irnW+WPKa7tFrq3IWU2ew6I39fpuou4jG/QBEHyG3tOmPZhteEk4Hhb0f4pyogm0Sa9h4GMq195YwJtiNL2fwuQ+LsVfIRkdOsgMXPa5MdcUVse4DAV/AcLmKtQ
ZTZ7Dojf1+m6i7iMb9AEQRaRvOFrEKNjNpVvAi+x3SGD4c43ulkHlsjyVirTosgUSeor+1VsbbG5l68CKHhk0hUILneXtFO+h0anLQTjycMe07czZ2duKjmUJjU4wmLj
BoMiHPw5GySYp51IAbs4wcqIJtEmvYeBjKtfeWMCbYi1ae5gGLv4VOyVHTA5IhxdyAwuogtAtHOIvSnNzuZuk/7opcw7Vcxv79sGHTNEnQVCIf7qwLt9U+/9lG2X0qvj
nzkDdlVmwMM8pfVn6MP0k+8qO7Efg8m3NhvLTrNQxI3I/EG6CzJ/7w2hwaqqBDXcYE7I8HRdiomOjyQ2q1k0NBShIb6dG7tXeI88/Av5bQOxeB1aYBEhpzFZBeNRLDHJ
VqAzFeXECQd2j1TSNcEE6go8QwXtu5EP5GUZ1WADU425hmMZ5MGoMqgvTRXjzjOwKRHXipC/uTKgjBnRlOwMkB5r82wbhM/yWqlZiQ5lCHWFNxAS/jZw6A96qepz3j68
DbDBZXVA/XYHxKFmuNzdPd5poE47DEfT+hN/h+tRWR2zVn7RDpXjUiQzfTLZd1IrW+C5Elv5e65objnGA3sRO/w07NvtuqNA2rPAF11UX9admhbP8ulVJoD0NTG1OWEZ
NpTzaST8AOEDh8vNYaPJFZHbJ51Mh53PFBDlHP+czmJW5EPzpagrDRGy6BushIDupgXtC7GQUd8RP9PCHpwYBwCdOaNWWhjT13QwyMixRZmuHm2HJbKRjsY4/1WcRdW3
nzwvUjsEpzO6IAb1jllp3NhiNQzYvuy4sVLxmegsB8d78PjIYfo1Py8RU7HKBEHLnVIicgV0AwiKaOWZEHfVUi7TGzTJE5a3J0MaqQCnavO7QYp2Pv+BOtYgsSDDBtNq
CLAghKA2YaDVmvzKJLvAnVwyIZJgolqJEylinDKkvNSslUymHmIP2oMC6aOFQbjZgq8zCNh4hJeF3T1jKWc9AYYABjm14gAcho91quNd5vc+0ltDXCvh5L2UJU8oRhei
AJ05o1ZaGNPXdDDIyLFFmSka3cK0Mk2lCgA0U+EQ55XV2Qr+Kpi+6S7g7Vi1SXBQ/b/oFNLlWrujL8au0xGVPjPOUwJ2jvs8BlP5P+jNDe9Yry+5J1SUp0Wrrw9eiBps
47oGd9KUP/YQ0OuEl5zGRWQF/z46i85RppQFhS6Z/yvFD4U2EY+RwCG0ZuZMLYF49H5ojxdoFGD1KvFEAHlVCMkFuEdor1mp8IN82deyT7+NJKnGePQL8k/ZCy4im+m9
S6XhH46R7YF9vj8zSKNQX8p8MzZymID8RZcLzQN5g4K/ZmatZ8ol9dL39Yz/5ib2TgcGvJhD5IQo4hk9XQKZSepuNQBkJGIOvHhYkPCY/0WSaJeCYGYIMsZrVyCPLMIX
bCn4ciGSyWhk7pd1M8siQ0lQ1knTtBtp+rYDR9CWdKQFWoZYE1SKLIj7KPg34548nER/KIg1OMaNdNdyxVjBZ0REIBBTfr02frbp1OFM4TgQLsVeD52bCwE4xlGFrvd/
ecN0mDlyefLoZXGmNw5ulc15In3Rv3xIJGDSEqlMrMbwIxs9btbSw2+xLYfuXy8T7xmOVlHAxOQo/NV8oYNNSCD8xQp5q5HU3YEQKVZYAJBslIPfSx+/ru+b01000L0c
+UaZi5w/xQrMcnOMAGc9JwnNupFkxzGyV9G7du7kfdS6YdwrRH5h8D55kLfMMps6XavF0sqW5Da/OX3StwHf+N3FOT5SUqQEx734d90Ydtz32sYuM1PLz9SoqFe7w/mn
SqnZvkFKMUplJqtmfleTlgwWGyn1g17PPxP6Fqi9MRyEcpz/5A5Yue5UTw95h8AYK8XTl+svtnNyY1TU0YPGrX0Jcqk5kG/Ay8USG4IpePFAxSYJMCCusPtQrmkr/3cw
9ju1IOJ6uE8gv2LBiZk1V6hN/kHZfxJiD9HGpA8xqIN3uosvdYSqDZ3oWBbD46/5ONvxdC0VTpvZVw218MF1lhyTwAbU3sCo9/zwWfjqayFt/66SR1gN9B1+rVBiCnos
IoX2zg4hddaRjezQUrBfyB5KlGXRhyec6Hiu0N4FTFYft9GoA7VYnHqogM99dGrNr9/5jIYuhry0/E6nSgunF4mP6hIoQaccpBOA+3SVG0YwXUu3wCGF2K2A/PqYUUdc
/5GhYMQZij3MfJ0rkTCuhTUfzMzW47pi9tSDVHbyj1HukZ2OXGik0tXbAy/KG91NehYuK/jFvBzMneExse5uM1SwLVRkOX25vvUtbVi1nFzfEJcuSTtZSNP8GN9UHRP5
uBNC5f9HkzbIdn2Yst6+usp8MzZymID8RZcLzQN5g4J1NT2ys2xgOoynJuVlTVW8bY5dVPIMi50kxj8CrCcLXL6yWYVHC0c0nIqh8riQkhQh9FTusFksbamkU4xn5VFs
7RisCKWmxTWIB3z5VlXB8cp8MzZymID8RZcLzQN5g4KVX0FXgqb3I35CCg8ganSGiNvFr6YP25Dy9rm95GK/4sp8MzZymID8RZcLzQN5g4LRZTOrlV5KpNQxzuY1u4Sl
2X1Znon7651Dq7HB9+Ai+5oeilK6igH1Jd588E2cnRKXXOTU2YLXEImnDz5y14gcvrJZhUcLRzSciqHyuJCSFPr2pkaTdqs86oodg3qOu+tLYUM/CVra8f1Ea5Wpy0gl
QBr5hWNCEg3AzvysBkRMKy15jW5vrWiDsV5L44OQwPQ5wTtUBV6ba17IH48hlLk9Xg9nyrTG8LbBfMQqmAbK4mCWyMccRrxoR5nCAHnqouhLRkMEA4wwefRuukZwWJ46
teVfqy8XcNixAQQ3WCAyKb6bfAPQw4cNlTn0/zDsIIxsFrYVo3II1imb4fOmAP0TwzgFD4kAKQyVK6Z/Wp59lDzZqi1BE2LcUZhJKR3ZhlTNfPXCVAm4gjKIc+SsN2lH
xU6f9KWqlCpRd+Sw/Fe5Rfke85DWsINbKeEViANagkKaldS9bTTK3f7HX96zq4VdzWiIHkvoMQr4EicSCust6ETNQfKJpiX43VPf+DX856BdhwqvhvlzxdDZR+2O+i42
ak+rwp/NGYWiyD6H4TsYnll2bN97sK06S1u9wC7XadW8bRIziTY5PycbNW9c+JxSk/sHpAKzQgDiEXuekNvLoGJu4OJ43r/pgsYnaHd3zJKFHEjseXx6247STIxngcjX
Jg+NsR6oEsVEFQOQJCjNnNtknUGg17jm40blznn8JHxJWQWKzohLw5RoS4YLpSMAsWo3ErUybmAFNSfTIeBmOrlJn++I2nr34CUDxN/37bspd59TSdaKloYYavYbAPJd
2URRb3e/0U4myMd2rLFFyD5vroWCASKq7lwmQnT6S2wT8WA8nkIX2iF6pgpHIt3C96XTtE93To7mDSbGauZ/gPyWSteRgcH37Ypwt2pydD3mAX7Z22BPts5MH5ZFO0wo
FDt9EwHeU07K071yAGcHLYj+41bml+OhWPwdisz+wZqv/bAU+Zo4QLeGhP/7FeBAewbiPTO+zy/tubmdEWu8JclEzf+SXIsgY82+KlZ1ejvOr/Iz4X6MhnDDgxZJwPUU
k4wNnBj8zWu/HNNYuUCiEXavGlgdP9+kT2RP2l4b541VpO4Dc/uXm4KlvWFNAG10AcTvF8gwooMKmKArv5m08LeDLIjYbYF9gqGKlRJQKf69wBV3afOpeul5rv/MCUgg
qjJqYyDySnealSXY4HKV/vel07RPd06O5g0mxmrmf4AhdXdiKJPuortVpF6gsT0uFmwNzLH74SDH8apHMa9lx6H77O/ljoiKpdvB449yheucnp2MTYHQFXqxWeI0VzNF
GeHV4TLmeO3FvGDDcNwf2oU/8yJUbw5ONaHM8eqR3ac7PhXKMByD1mWP5zAXAUNegQb0GoFcxJTvlLbu3HiDLBCJLOS+HkbD+vejgUAUYcEo+rsZyDPT061ogHbiPnN+
RqzYxDQT+5tvVznLzRqpK6Qs441ylWYO/gVnXw/scRdAOycLx40EyzLtRpAk+ct8t50h3YbP+u9syWuxY4+VmpUl2fJT8Ot7wRMN2b+G/5tOSp2/7M7gQnLflX6wqUxI
DaCxRn5y2rEHEv9pMyZqiyx6+Vyw1KYn91eWBz/exQHG7xWBEWDXZNQFTaJZA6/pqNZyg5NDRhN/VY2LPtVYefP29IbAQsfWHuNZ9WYFNqkoyKarooTYxVC91FzejkRv
YM19dYvShFdh13e+CmA7OTYAe7uyhCvTRMMOhfjN2dRSx6JXmw12yJXcZz+bIQTVsdPapSbSq+ndlDHuZYzX7/ifYfiqLxgTAmEGvzI+TvexX3v5/ATtDgpllwZaz4C9
DaCxRn5y2rEHEv9pMyZqi7xV9r6a7EmuVY8+GRGzi1isLw7kDWzvN0pQ781dqsY9313YVEpOigmkFXOCalIhxe06doUuHTcENhrmzqomGWQ8YNTBkX6d+DST6ljdLj1Y
gSEUBihJp7fQjaAWxz1C8lJvuUesOQFMMa5T5dbDGngIzY8WUmwy5FiGK9hPwvI4UedDkQMKEp+HsNMtqNLvn0SOKREwPnYsrHt9s1X1Fk1RovCvkF0Pm9LnK6U/f57T
sTm07NUwEoEkkVHRGRuB6a7IJwfc0o2Lng6NZiBdODkLRF/TRruBvOqD0D7akIFRUMTS8TAReh4bTegy1voU302lQqtKjAJQ39ITj//fC89Oez7j+D0tlR8n1bV6wYjs
kjGe3LeUdd0XW1JxW7At8+/rmTtIEyEm7LoPST61DmSSbnhdbHhGXv4n5OEMJAmnUa+e26Ytsx+XdC69MzF3e5GEaf0b7dUecROFM3QyNIfmh8lFIeRxDLOamAKWDXwB
lWeZMokTJIg6AFoX4HSGaQkLNnCTIXJkvthWC2W8oa9NpUKrSowCUN/SE4//3wvP5EO9KukrlxaHIpWujumltFGi8K+QXQ+b0ucrpT9/ntPrNLH/8eL0dzgWkcGkDUve
LHkS36RkAd6XqiunGV08+c21e3uNNctjXEmUDsIaJ1bQQGpAT/4GzzVpmDbjO6Yk/CnnPxqqQiIpsMp50VNtB24+QwcVYJFl+6eEDtgSp0rXbl/rxMYjHTIJyM4Mqf77
djdRq/CsubYAa8eqmqos0P5B5a50rrT2HYcR2UMDQUuF5vh9stebumdiPKJAM777lWeZMokTJIg6AFoX4HSGaQkLNnCTIXJkvthWC2W8oa8f+pwdTMakOqvShf9pwAzc
/KOw+ZwENEpRCzYwecOfpkdsTxHSMe8UaREA9s/I8YGpLGhB9AXuNkuaXiicrj/byogm0Sa9h4GMq195YwJtiGfWk5t7SYxhWWKXGkdew+4qQdNgtnd4VWBHoVyrxvys
g4vf17ou6TFWsb2vPLfYsN7YN+iWSI0zfA+1UPUf1bJSmokjgc5A0+0B6JqbN9Qt57iCF+H4/bQYRT4K7g2F98Zc0RIJdleFrDO3f57S/BWdFBHf9cV3apcg8UjLItQN
mzx7yI4iBEQiSNRh+QT+e+drmd9h9+kvGwRZyYKC1CbtkNU9raWPVNCHn1RbVn+1lHBEs381QoTzd3jX0UKdfMC9p02lfpmgjvk9xmVcYGRqZpLUjGfSr+U33lQHMLYn
ZH5cvD1I519gISTuQsfUGzmRrqzYXhIZENtNRSzRe8wONv1dK7UVr5odHHDk9HIe8VivB8BhJIJlrYH7AJkVP/nPuR/xWN7I8qPFFdL0SlerjJ67NU5dhaIY0Ejh3POE
te8smoFFfd9RkC/BRMDxBR4XPFM0sAl66G6FvHKSHcFV9PMZ4TqyMzpoQRaFxOuDAV4GiD20b0eDvR3T3iXj/yeO6ZdjC9F0rT9N8lvp+UnLcCluFgQ/eavJPCjVnsDA
lQu3QtL4cc17v91ef5tDxzPkxWXkbEZcuk0UQ48PJqeOViNeqoUSNEWZBRRSY/lBHL75EhoHB5eW5vXYt9vzDItlG5Ew0kEi1HUSNFn6amS4qrQZDcwWujDcuwR+FUoV
yUCV13NJlfV1nN5KRnudHsxjUWUzqmPXw9o8L1XfS8/FKdabDxKp92iNJg/MbI/4CZvM8TFuFCkCBNGL9KqPIDvK3ZxSWHO20yonVBuSEz+kOQM0e8u43c/bte5TKAF5
JkE3FXvB0wVZjEObIUlyWBftRiG8YZmUJLEWVEmyy/VtdeNJmncnuUi7vCpaw1xqDE46wI9gMzeHnCuT/cJzw7lJn++I2nr34CUDxN/37bvXfwmavFUpEoZQfYCyzAS6
pujQJsyEfGPMV+Oxs/IC+Q6cw183zTzpIqYbNQjhG2YpKuStZjZ0In/PQ8+nS2TCSFvdAPpxVKQrsD3NUaqo57Hn2KsGlmp1whiAV741HlexeB1aYBEhpzFZBeNRLDHJ
tsldZ4jcP5npew4AGSvCMSrt6kELSYuU45P5N4tFqV4lIDST3vyCCBmUgy0xvvPqcxiPTSk0RQLsCxwbfLWjJLbJXWeI3D+Z6XsOABkrwjESGxlgELeoV7mf/hcU/Awj
4TFgNp2mJ+AOUsOS6hfIOge2mJI6+aj1WseH8cO0AR4PS8GSnHj4tkfhTn2m6ikiTHRTzhbwvzHwc4G0nv5ohAh8QdlZyd3MKp8oYsf8gCC3V1B01CYIgzD56oxLA1bm
2zE0GSJPzwcDdnRslZ0vfBEkNYbGy276uH5T+bexoYCeirM/AcJydA5OOxgCMFodUnUA3y6KEywOdoaDLiqkoTqpuJnGcVuziWZOVWsTEiEamHkoCG+uxmLRohe/Of96
0MSPzr3MXmswE6n9jmqm0/Msm6nfH/Zn7GN3LKatcQR5TCe09TSHMDFh4f1JrkDi1HKBntvrFOHd4shnM0xsUPI0AuqMO2b1zuYLl77NnQFyRKxIikrp65jCeAMKHDtJ
WMqxZfYNCVYPQlWQjcfGXRn/wxWElJHHjYq7i9XTW8ccvvkSGgcHl5bm9di32/MMDPu6yTxRjR03fEqnT06nGaTMKUIahdta0zbRNsLGyIBlzgfYY5nirH9J9NIGwHHK
81V1Mw8u4NMgjprF4apt3zAH322Rgt5d6gSX0CRXjMpx6X19xwaGlw0kVZ9MLjI6taUN4R4NZu/jBZa3dK9YRYNnrdy9tl9eQLB9SKlfksHK2TSJfSmSATH+1vmXoOU+
6b4vaFjMPSBDE3NIUNnXKQmiAinLDIWWbmtE/DwijdV36TrLUyFSXwSQPEGU2mtz6INE47i8Ol/YJRHFlHfwj6cAL4mXyjRZtpv5u/3ytnZboAymhAFDPuqXJ8FxyvMK
8ysDNvmPpUDmZNqAt6794AWwu0aNhzhm5fvqvqIb7mC3V1B01CYIgzD56oxLA1bmM6+CzVWE5izLSMO/1Fb0/eiSV+zzZ0H5tGg1DnOSqHtD1GlsFOJHnLJa47mD5AeD
2U+Uz+4fvQL7VRqq3pGzw01joPcfJekPDP48+LuAgVn/wZFbx6x2GM7wsZ9LgDHVub8ag2dmTC2EFWJgVnd0VPGE8KMO7/WTcQsECMSWi4CrltP+f3woE4FS78aFyp1P
PIx2HHI0rtcreYuBN6ZqSyxCp7SRAvwz1tYMc5sD7Z6lOhihgwOCTy7QN3cvq2cgkLwUlNaaX0Vw8C7WPg2v48DoVErTNtMR1sfZnneGpW82q8LnCgh/iup7IrcLpSBl
fF98oF6dOtqD734DYelBTNuvg9omMitogCqRQDagHrgNLAEzriM0jyKYzcf0G2ZTf2n4bjoj8COkR+Rhnnzh9MADsuY7davUFwXKaQEum4ooErNfhNKnwchbJB5jyUa6
nX3rkuLC4L7kz7agLTDNrvr4GXkMRdi+FHpW4Ac061HYancBmYhpebzTE3ulOqwLBDS4KpYUMsXgYZ66V0uCdSgkfX3Plnk62ATqrQaSU2r9lQMvihlcA2gqxa4WcZjL
6U/+IESQSj23l85yNz/8N1MIxluwNKM+3c/ewjYhDY/Akk8sMWgc6G3xoI3RoCXHD+wG57oTFLCSqoy3oTNxVJpDgxWs+SPaWsDOXm3buL2lPDWrG2XP032dE2YAKwyd
Vz9LRgtpeK5TPAO7nfpMj05yh+uOxBBTcQ2dpKkolom6jQqtY2qNS/gbwRaiT4cbVfTzGeE6sjM6aEEWhcTrgwFeBog9tG9Hg70d094l4/+b0t5K+knF+bhDXasHdw+0
jLU7ahixfCmerYwW9iDZ6AOh+xc2H09AugNP15uqAh91krnWkmeEYkFVxOIyB567bj5DBxVgkWX7p4QO2BKnSmCQfr3CRHFKjQ1cZdb0WccbNFFRFLKq+gqqjtGzylhJ
DWnRkIWi2piUBSYJVs2ODlK3BJgpWT/bhvqrFVsWdpu6IxmzFxzXk0Gk+zU0CX0NTsUOyD5niTV7dzvmxczSk+EJ+s9D/Z7T1zjitiMVW2zVMyIL878WNcaWxy14XY0K
yKyqQfN5nEnO1qpIAlmEbP47KYvWPQU1ci5BZQwZemZojGS9UnVnk47i/9McmYmYDWRxR7s8y5x++9P2iJyVftb7I+NWMRKXdwveUlUURln+7yWlPHloFjgYtpga3Lq9
AQFgpan8T9YT0aRRARjQ2D0LoX08b6uLt6XGCiBpzpyzHCIaKJNsqrnEiP70soe3syBQhSlve6pJsi/JwvrdMQYXwmrWA7hOHEFU0y681qKkLZYL6uR6f2MDl/DROfp5
/bGOAFRq6L5eqO2CNnRoYpoNJHxjHZQC773lDRMBQOGGBAXa80Ou5uaDoILVmGzIZI2+6MJGwutF71SRzls8lMYxYYnpBbY21OsKIXB6uJS6/S6bHdZEQeiBxkleunkb
bmm2KJRatMioOVi+uuW9zPxrW4MJ/2Y5r3FoqvE296c7PhXKMByD1mWP5zAXAUNeBEPxcLiNr2uGwvhboSJH76KycSzwJlSC5w6ZXLxK8t/B51hOD63lnzcz5x7X2MCu
1xQpONtnWsNvijx5cvFdwICmNxzirTYd7fXcs4sXVIRYBfRpKryN0+d9ih+DdagdDHaQoE6p2DKoYqEYo51/TtkEJWv1V8aH8oY9VMasQz1AnLHmwpJ+Y4kojhtHL3GV
9y1+pBZM34DPxuszd7oMtqLNv/rOC2VRacSIU3LCmLoKMBqPH9hiLmOpCENlLqVwt1ZVf1l8msCL2iFoh3pKR01sCCwH2fCpjUATDI3nT+c1K76Ha/tLSgr2aD3/B2Zj
I/jooot0bvq+VVQM49CuILMHHqgXeDwg0iAodVpftk/TFl8kln0OoMsxn6Cl5A1DGxFuD4YDAur8cWd2K9OLYr1kVCqlYRYZC07/5l5IFE5GsBVRk+W6u8jqxMIkx7Ge
qhkZNjShOeiUisSn+Hj0GvVGSS72NNeWLSqIPBvh4T5vZz8WHCAWbvpxrKsuEkA/ItULc618HXW0v20ATT56R5NN33Oj2BdpzaKaV9WGQv18hz4sViIAFjhlAXnPznmY
ho0xuO3KhE5XEEZDCVsr4t73PWqsTBnhaWhDWcrifYAsGonh/WlzTvAzRlMQ6JquXGzlseW1D25zLj3FDX8HNmPimyZJR/F9W9o3plNNX5GySPEYGDQSfRfobLUgRkWH
5yH7G10FFC1zNWcVIDN0k7qE9irs7nRRh0AKGWWSevfV4sLom+G23LtYl9EzE/5kcJ5HPLnLTumc8oWfVF+UQY/m+CTyK1uIXUUyFuccmJ5uiqyZR4c20sSPg9f0Nn3e
xXZaPpbyu0QNfRP3tkbxFD/aqxE+nhezx+L6LFdldSfo5NV2cTYXIOKLO1kSET26UOFJwZAyKwEwZu7HtI6lfHUp1SuOMh2sQEue9GtwC9sCxC9XtFYWwAXUc/2obhMx
TGJI0xCXYLvLtSc0EnnhCLz8MYDGRqjjMivYGuJ1H2pwnkc8uctO6ZzyhZ9UX5RBGxFuD4YDAur8cWd2K9OLYsAFbbMh+7gGgcPcRriXyTNGsBVRk+W6u8jqxMIkx7Ge
lVhRGiMbal4Cu8Al5BytbFcTdRTMEVPD/QSGv1wLnl3e9z1qrEwZ4WloQ1nK4n2An3DKLUVZd1Rpacl+2178/HhCE9Zy7kzJmZxfRn481SMuYpGIjaUi7tf3s84xauPr
+1ZgaDg5+uhuAP7eSrzyylDhScGQMisBMGbux7SOpXwcTq3V1MatJieCvrOwe9mLa9ZPeR80K3JGCHLz5NVAalDhScGQMisBMGbux7SOpXwYkIqFVY+pYCxjgqlXBb2o
Cjqe27PCcvUhNrC7eXBOhqROmJnmSMsXMDBbPW2w4O99waJRCfwZ1vGTMGuwUfvtWOzgUHHkNI7QjHY0wAqiRZyibqUkVJKJjtnjdDVYDx2DDAbwQOTsKXkBP4PE5Yao
HKDSoxg5Ue+FxGQd6ymJbKKHpbFxny5DovaT2BmrkSzijJr3D21a9bgoc/xko+/y8MP2BP6E8PiXN6yA11NutrP2046V0iQ0tP8vEApaipJxWv9sHrRGtt9/zw9mhZkX
I/jooot0bvq+VVQM49CuILybdr2dLZ22TWL/829Pon9Y7OBQceQ0jtCMdjTACqJFGl3rYtXhb5gnMCWuttfd5Dx2StaJIPmd2GBd9Y4jCwvxUTun3TZ83cNOIjv5XezU
i/QnOz8gxOJ6k4GYw8j+kBdt12PBKYjBrtdScumn+Zub2BNh55TQk+b8gwIF7NFpMcDcrS/rGEq01gip2YmxVr1kVCqlYRYZC07/5l5IFE4rRQPV9SFNuPBfOqrVkV3m
P1gDmwJmD1qmgbe1YadBdcqIJtEmvYeBjKtfeWMCbYiPSmr/yc3nKU7PkMPB69f2h1a5EfkWPkuRlUlaFKeQEKgIhbAcDIAbaGkZt2LREVMlf1C57VA2vFbqS7dR9t9a
hlRyntLZVu35OWoBZ1JenQoGwkM1er/PgcW6/yWpSs6u6X+eM5v9qUUC7aci69Ud+8YmrMsxj/OW1BVPaFck557vSXniLe69mVBGAmZASRD4njDMv+Fx9ewr7PfXSi0u
m+4BpnkInVGc71MgMa+s7dGsoZ5dlxR5G17tWX0nfPax7IyDPM+AVhskJSLMfSm8Lz8izTcqbRMp3QJcpRkTXc70JIKg4AtjTp+uJ5VBcY3FwfsqwZ1Ii63z2Nxe+ekW
HkjmOFDpIVuJA0XXXMjkDz+WUosUH1vyXUNjD0pN40FQI10OdZ3/iyvnAVFVsTKR1AYlBd+Xs3VKgnjZ8WsK/bzTWpBvK1q/sPeV0Jmj3pbrrgqlS+ZzL8o4A5Ia4eX6
KlbvoBPNRUZX4FcODJke8Och+xtdBRQtczVnFSAzdJPVFx7xVeomhTT47fBmTMFUqhkZNjShOeiUisSn+Hj0GhnCeLBoefiMUnTgjE48OJ1ZpsJKvUxPy2tT9FysdP/W
3zt4axfqBiS9pwGP0e91kWv+fIUGJdwAjkHDepExcf5Sibb1Z/giBPe0UMoruFZcb2ohrU9MSNQ4fdHW7AZcl9QGJQXfl7N1SoJ42fFrCv3j+ebu/uJ49LrADT3VvUVj
AqwS6KeiNHCe29RqWW9F/wbVQoaCqpI7stQfFyd5gQrf3Q75q1kdZ0VW6H+KDUXM7Qto4nWMnEGhI2nH58PKBJe2d4mIOHexA+4XQcUcs/dvURZjx4/SNbMeq6DfXOlY
hD5pzYkjVUKN3/2cRxkmBBwpACG5YtG38HqqHpXEnXmXMCDc25OiN1PjAaUxfcOb1W8cC1ElOejq4eSABeGCnZcwINzbk6I3U+MBpTF9w5sOaOpNxnYMeZtu2s4EcG90
7Qto4nWMnEGhI2nH58PKBAaMrZyQJZIQFGiR71ov40aR5X1Gvc0/iy+gUfVnQ7+sYL3vMpjZA/eO2aDmjv68BcVhaxZAqpY5Gh3Gx7wBjVp7Q4C4VDw81f11j26rH00w
iO0jt42+QldAJEYy2gjsNct/H4NH/wbjjVE+e3c+RthE29D3JHGskxIUD2MWuBHwLSfUOgoh3ryVK6DUxE0hpUzEfw3Spi7kcPDEg2tYzbcbK5SpVQbYljOiVnEYVBzq
QsM/IrglHuKaGjh70qT/eNRZ9LmkTuXk4ZTMccZ2Zq5Sibb1Z/giBPe0UMoruFZcKQEUuZZ7gwYlXWtSPvg97aKHpbFxny5DovaT2BmrkSxi2RIWkdaZQ830XyjwA3sq
fFIGyzV9maSjgiFARuUpId87eGsX6gYkvacBj9HvdZE8PtIDHHoA+MPE6d2rZh9IRNvQ9yRxrJMSFA9jFrgR8BO63XaKILQfaBv/Bywku6eR5X1Gvc0/iy+gUfVnQ7+s
4oya9w9tWvW4KHP8ZKPv8t7i2i0i5vDTpPKhVKSsKoW7mzkS3og1g1UH8BSLEXfEdS7rhI4kT5ucgDA92PRYpihjCialeFGfuGCGETt6jASPeKL92PxpFY+ZikzYhF2f
e6erSMhMdwmRM9z0wDyx4xsRbg+GAwLq/HFndivTi2KClYaabgh92mQOaX9SPnisGxFuD4YDAur8cWd2K9OLYv3EsPnRStfs33S4TGRDQq+7mzkS3og1g1UH8BSLEXfE
nzbPyZzjG+j+J8hDVK7FTm9RFmPHj9I1sx6roN9c6VjIyS2M9Yp2YfSPs3zSsS3+imXHwpRak6ScwGsZp4uEuxaZMMdmcIx3umcK8L0g9DZC3n/GHIQdAm4qamRyJRSE
DP1sphVyYv4n95Sk6Yp3OGVNgyZRjvkHRNOT6Ylizqp7Je21t6Eqi4DqyPYjCpFasP5FMcZjR/hkkF2vfnugMTKVI40OtFdp15GOTDduO5Ff4XPT1wOTTbLonIgLwxg9
MD1zfLVXxW13yByHnBevSUcMDgwRQnErUzM0dTYJBThc87IOTcgLSaToZt+lYHjUzEmc634dxTWmEDIprOIYo6Qtlgvq5Hp/YwOX8NE5+nlfk8o7yC0bDaTdHKWeaL4l
WZXfHiYtW8E8iW8MhpiSB7IzLKgpIq7y/jOqPj6z1aNfxD2QS7EmhakcnXZAOxCHUC3Vmu6/hWlN2nLFHqFWj2Ju4OJ43r/pgsYnaHd3zJL6wA+UNgMi8Z7Fd2/CWeCT
5YulsJuxllqZGn0v6sEgA9h7GwGnxvXVlBIS0QcXQJqv5q28iLCdplkzZxNtizbZuewhXLEBzkFyeQrd/WsWHeY9wofYoU0er6HUrtwhnRrUgcyDVvDwzjtIkqkGkLWp
iMcwwZHv1D60WennswBHVKrn27OIyDUpFM18GbiQ1bx0m4EEG9mVJ17dWE5OAOZ/wZ47msNGujOSIC1pleQzEyft8njzoLZfJkjVEA3GUoodDzvCjNT77i2NpjkAPOm8
JOyEUl4iRWp2vi6bYupMwZvYE2HnlNCT5vyDAgXs0Wl552et238vJqaJkbGMsJgFPFJqEAYjqFs6oHO3seZLQJvYE2HnlNCT5vyDAgXs0Wn0mi+gZHkZdo3fV8ANzOGP
AsQvV7RWFsAF1HP9qG4TMUYTycwva/p0eVy8BgRwDGzS39wPAxTAkKHH5V/BN+gf7O2xYwkn9H4pHbQwPc2710LDPyK4JR7imho4e9Kk/3hjRiGeRZMxqBXBd/ooD2Ty
wBzToZTWGP1y/HEvRxdUin1/RLNCCHDHhFMuJu7/ikauFlaQogQ1pN80R6NVOaum0Crq5hsnlOJsVJMAI3motrW4d4aXjSq+l+HzDkFvRj0vfBgKPkl/IPTbg+FCpf08
4iodqyrpkK5ghLDsNI3s7oW+zQVDCQI+Vp5L1FXFLj2rCiFnGo5t4jfLT/X/BAsxUom29Wf4IgT3tFDKK7hWXH8j8p+UyDkmlhSueoDNYJjetHwYEpsMgmn68372oz2V
fX9Es0IIcMeEUy4m7v+KRql56hFsdUcGWbuHKiLMwDfK77RB6IEtqVOQ2ENBHstx2OQFJmi+WpHEvJJYCXSZC4YAlGNRYn/OWth7FvEnEXY9WsE5yHem6lFRybcPj8B4
2RSRGFSm7XHFhiZdlmAk7bZMmcF5imb9aMI0jpRxg38a4GA5CQIF7eHEJZNf2pVtiydldj7wohBhDviqq1KbUNnjT8zT21f8+t/ID0HfNj34n2H4qi8YEwJhBr8yPk73
4d5dSVqsfq96K+mZGT+YPZADXdTtU7/HobPzQUNUUB97k2x/lZfmsSlOaWtBaMX58qq4+U877dEo2Sf7T1wazlKJtvVn+CIE97RQyiu4VlzFXsZZIzYcWW8jfy674uEW
wedYTg+t5Z83M+ce19jArqzeFI/xdVjQL6X/HU4Eng6xkdubgOAyfgyIxZC5MrTFUQBGXQgZOpOJVE9bMGqbO1o5atVqlH38iDZayGtY00p+skbKZhLr0OZBycpNQs/C
tWtHCQAgMoQr42sPKIcpFsrvtEHogS2pU5DYQ0Eey3HKgYAmA+nW+CjEafmwnGcg0QvbB280v9M5XJDK59TMDoGtQPQJ2wLRTcjuy4umckRgrL3bOrjUJ91cgceBjQiL
NVL/vhZxt46hbH60KCssP7k8OsKRDE09acnn9hwect6KN2VpvMrgxGAg3TTfmvsFa75nwtG0rWSl5q1RoaWKWH6yRspmEuvQ5kHJyk1Cz8JS91hQKYMUxip5sO+MhK18
yiLwlfMt2Yivn5shr19z08YxbeozPejBJ4gDsuqOHR6XMCDc25OiN1PjAaUxfcObe7Hv6Il5kOssjJKf9XOcp2uOQEBPgr0W7RC39cz56aLgo+9e0FA1pL9IC6EKpod8
DaCxRn5y2rEHEv9pMyZqixgAIbjNjYvaH8g302shjy7ItVlA3/sRQe+PaLvyCQJzXO7hHnk/duC2aVOtdfWehgQxr769CbrSfk57i6sxXHOolGVKtK/6ceVvqkGCMmBV
OnOJmjmyJnrMdW16IoVo0qnYPxEvX4GdsxAVqgVIrYCwv6XmLGaU/dbkr6ra9uJn+yOy1JByOyaetKeuBcm5pq6jnqOGVg3gN/TDlX2OQidz85KGOCdgMGccuMhJHaqR
AR5S6jMxPzN3BAUuHt4EOgCZl2jyncSYqF+/87pgiYtQ4UnBkDIrATBm7se0jqV8MZtpmi+hpaWIkYFOadXxZSpyDAfSnH2R1flpgIjDhkEQiSzkvh5Gw/r3o4FAFGHB
DHaQoE6p2DKoYqEYo51/TtoLIuHJNv83FZSdsEeH3T5Q4UnBkDIrATBm7se0jqV80OZX6XWc4jbzoVY649zGt6l56hFsdUcGWbuHKiLMwDfEmBPSk0KCZ5KTVBLjAZeB
eOrlEqKdGKAqDcSRP2GkN92cUX+kBd2DoV0AjK3UdL0QiSzkvh5Gw/r3o4FAFGHBYrydlgFKrbIr7fvsr7RDg7saQdlcMukZp24yAyW4DK6o8HDwIuByDKtF2VzeAPa6
dWYsC8ZMyy5lUfX2AAnJgWuOQEBPgr0W7RC39cz56aJCPLMpjaUdj3z2PpWhc+hp2RSRGFSm7XHFhiZdlmAk7bDiuASg0dtTcepy4T516lC+pqxXNZTuTjti64mtXW6d
1vQXo8atUjTrysugQklr/iDhuFtWhU1HyXn62aH2pxavosaY5QPTOMQUnCN7H9y5Pa7mGTRCmDXZ2Xf5OUFvde9irr3KyqisAxVH3C7+/Wmu1gRYdaR43KfRuRezx2A+
lF4OnuK8HPFlrgEpx5VfAFKGkgeD8AilntWFQnuGTDcwQLIN6JRkhWKv53Nm9rtj4h49K08aGem0bm/AE6/r5ojdH0Ii8RGMjGSbLQgTulA21edd5XN/3hBGKeSz/jQR
RmwRtp3QhbPhlnhkShslW1PwOFf40lQ2LzLJqN8XWhRcO5MxTDJ3OMEe5DkWWUkiqFA7xb78FJ+Kfq+4SFiRDsdEmSA6YDqaAFQBcTFWuSQ3VCnw3Z/8XY447nhSu0WA
Bbs5D3cYKnEqxgH48+ey2ypB02C2d3hVYEehXKvG/KwDySQHmRpstNABadSkweGyYv2IOFTjVCG394EsATiik/fMKBTbK9p3I2KKdx/ji6EGe/tgENTN+LB0m0vzp7QD
aFFfJxBW8+hVimc3Qwykrktt/usDp8EXCVKgYH+sbZLymi5BdW65HhPxBozOQ7bCG9PaC31nHDXhnskJxG5gdswKhUcDxqHSUenB5jK8Sr5Lbf7rA6fBFwlSoGB/rG2S
8kgeaGkF2IsJkmuSH1MWrtHpLK0jKzicihlhKeIfAG4xr3K4GjXI102N+opq94Dxys2gN+30hJi7nMsAvrd2qajHhqxz0QRZ8hnroNughguugAowZ86NrvytCrh9Rjuj
6oMhXnMmd6o+5bKNErCVOiO0zINw4kJ9oJ/830E7uhVEuSJHdAi8jw0E4/qOivzxNDsmzRCgJHdtQAkqwgcXmXKcYyBpkZ4E764l/igB7JEEtpAgYOL0Lo76R6BNJKip
4hM2GnkvyLzTclhTEwLt7eIBStD/iUhdaDN8iYLJDHEGxYafgGallDjuU0acebxcHx149SDrhJrHLhbOn7ieAS7alsojy7JW8maGG3jL6AMjPlTJc+aE7PSzruqztFxm
H0RBYdEazxt5S0Wj2Fieb+A0DGJAbPFvcSuKDjDji1XWvx49AH/PX0wm1B49D4f6t2YfnFuJiNfBUOB9CHtei85qrqxX8M1tO00SeQX42Bir75/pYtG2P8mfOQOQ5RWZ
zm4WMPF+Kaup1Ga0UEFZgduNDwfC40j+Nd3ZWk95g1f3HpB5cKRxuAj+OI3QqrMVEy1pzCL1LvT+jqkVeOFs4EjM5MdhteIjEvHWNW8nQNii2LFN9c11kTf6dE1Tdsur
H7qsns+3drobOr+zOqQIW4CmNxzirTYd7fXcs4sXVIRWfKxwfKKsLJ5LiAUvTwezv67pIIoa8T91YATxBeSVCKEQ+9crz1O5r7VOqCJq2GFX4RfFDQJ2Htq5GephDZXP
5yH7G10FFC1zNWcVIDN0ky4ipy5fuWQpLbi730eSBGzboZTa1ImTAJOLESKvBDJ6zXeVjc6XrfgOO3RQTAZU4Wgk3AzePgbDfBZ7qUDlSiSlefnFOMS/j+/pfhAlkSrH
3BYAA3Nu0BMXtZ60286uGrAtBEip6VSIMzNxJj9Au4SP5vgk8itbiF1FMhbnHJie/xnThDIgbfp5C79QG220G/Ya6U8DDDYR4G6mwpnCL4/F9Yt1WhkvtjuFwhdOJzat
g2liz5IxWJTLJYPFevMJmoYAlGNRYn/OWth7FvEnEXamLvyBFy0CDgiS43EwyFqXfrJGymYS69DmQcnKTULPwq8tM9P8JHKuYCRgwkgqj5Qcbs+bT8M1RLteiMzks48t
qceisWFog6KgshXv6CZ0caL8rMamPpUrP3AmOY436sN9f0SzQghwx4RTLibu/4pGhCCSQ44XSstTrc6ody97c6zeFI/xdVjQL6X/HU4Eng7R7RMI+0jihq7aIhZD+06+
rFvTQ7UNsu6xZXHZIDyxE4AFj8rF4B9pHrI3dK11K+IMx8sGvND6z3bFZfkwUu7wL3DTorJQgL79sAtJaZwEnBsRbg+GAwLq/HFndivTi2JADtRBjowU9FB4+FsPUrIH
Gl3rYtXhb5gnMCWuttfd5O+5QvU3X/yB4+e81zgcyLNRFDuaW2Lw0j+0uiFZSumMJ/aCBFfFHdHI184eyPHbzYNpYs+SMViUyyWDxXrzCZqGAJRjUWJ/zlrYexbxJxF2
GiEE7vcvT0t0M3TQ8OZaaIWgy2tRYn2tnqV5FJLEGa0bEnAOhRhLthJTOByZNhyr5JEdn4e7bBRK7kXe7K4jhtqGi2+F6J81iYePv44cidjrp2BTlXIIVt5lSAG4/Rh3
c0pZ0LO262TivAipfaG9y2RuLNACROes3dH34j8A+ciXHx9cgPiW+2bXPYwVAPPM1jtyxE+iAF/HhDWezzDiiFTaPuQHginwHRd0ZlK7P0757ZmHoDhhsLbbX9TcjZYV
O274smv6kiaTpm2eJyCIX3PyC/M6nUUbNd0QDHQHF/stkmJGjkDfTyRAtQXEUfGhHjpp0LWScdkpU0+e5tWbdJyYy3bVjsF0uU+Zjlb7Jw6KZcfClFqTpJzAaxmni4S7
Fpkwx2ZwjHe6ZwrwvSD0NkLef8YchB0CbipqZHIlFIQM/WymFXJi/if3lKTpinc4tjC4W4t1o2iGvW/9MyPSVieWbhpy2UFP+qfu4YLKoiLKcAFy5/BwO+MriOkUGoq4
OSxcStIup3SVCgDO5Wrceye7xkFivcbDCIkOWzxtlY6QjvF0y0pr21G78pP8ytf1MvIvlKNTfYYMA60dFVIJcDmwccfMB9FLrafTALGAt35b/x4cYluGxqHlxKXZ3Spf
qu1ZBNs7VjCIne8KPL777/ldgBLfz6DZHagUwHWa/qzb9sq2WyEAh2N8vJ26EW1GUgy6Jr+RZMNVbfsOyO5uaaQtlgvq5Hp/YwOX8NE5+nkAcmBid61FsUikVpKpE1wa
jXME+RMUZidKNgjPXTJrUIzBkSc5QeW06985u5RToqokr89gK0klnKK4vGahFHsYMu+aabPCZXQQIOPryomF+o8xza4Zj/23AcEOs4yCYwGWcK1hDkSFOwlCwCTtZVco
7ido+ZH79zRJzpEouq5daKbX3c5EIsgdTiozNBoniqZ9U9DskQHuxxaK10u/uU8dVKMlqXSp7xUzZUkO/dbS7rQpTBn5f+Y/OSqb2QS80Wp8KEZgIoBeZwUvHa2AfIry
nmFo83c8IazQxWNbcd6dvP+AaQYKKgNcesR8URZ+aWr4n2H4qi8YEwJhBr8yPk73F4aaoN8MxPRvcQgnyt5c+JvNtUbl4bU48pW7HnagecbS39wPAxTAkKHH5V/BN+gf
os2/+s4LZVFpxIhTcsKYuksEdLwEm3SswL1wpbERHA1k58NvRg5mXKM7i7uZVmc2sgIttEInUCpKFAodcmF3YBrgYDkJAgXt4cQlk1/alW2LJ2V2PvCiEGEO+KqrUptQ
gThzbjUSiENZ9YjZ+gdGu4BSodBNruHbUYfqWfkt3t6W7xXDd0TbgIv0HI05FaM9HhTCt82yE73VmU8ppW9+PutB1NGMUIgCr9acgOS9sf2pXs3Yp3GucCMDP1s25ofy
n/hpH2IiGpTMsGN8lhPt76BHQDfW9wnDZDYozwtFJ2QdDzvCjNT77i2NpjkAPOm8p91rsTzRsuT1HqqXqC9uuD4jTNY+UwdZJkxFZhFnbTh3a9uu0DcyfIwTeRgzsjpb
AZZ76U1pF2ghA3rc6ewOU0h8kvAjfSpsqO5fPrzkez8qQdNgtnd4VWBHoVyrxvysWYM0BU5aINp4uTGkC0KnUZYU2W9YYbwu0Xas8wC1/WDYd5iIXkMvguaNk1JCYBwa
5QWPJ48i3LNmcn1nVa3RALeLaJ2f7j7IBdYIP23B/KspGUiSWR55+Hum653XZEDHcu95DYYfNymeqa4VlTybAFnAW5B0cl8vkLm/pOAi5YPPIch1nSogdziBCFIacYkE
k5kBlDLA4y2Li06VJXX/rP18JA8ZcU0XwL/seYS6Ea+/gyudc9JxOQX/+vXtdSklB92wT3gF0trMVPS0iFAIRWX0WsCBV8mVQaRrdw8kNr1HbE8R0jHvFGkRAPbPyPGB
Ez4QP+I4c46n4nK9vdrMdiKIHEJ6fXFQOXJT2eN3jfQTTYAk3D5M0puRoeEy0SVJd7NeytWasSn0iiVXgB0rnX6rYwpGcr4E2Uxdh0mXvMakuQFx1sC49UO4a+uZi8gN
UfEOCaHxzdrwOlLa3Vj9DTlrf2hXCVN1zEJbu2INdUzYjHhL7H/Oj0tmv5uzFN0si8PcD3kr+a9XD29sOD7MP7pGPjWm9Td21xrd4STsflqjdPX165rjMppSizDyXGXt
nzQ5XVV8X2gPTlMUP0qaI4uvyyLDzmxyBIw6FYZPLLR/3re3cTkfgp46/VJ36OzyEz4QP+I4c46n4nK9vdrMdv2Ij5a9xfszgEzfbV7Q/fmo8rglXZLLyLc2wTo9UiTs
nFGmAB+mScq7/hceCGzvRPU3t/DwQEJCocP7+aapLRO2/jkVQsvTzPbbjK8gyrqDqhmo6irnW+WPKa7tFrq3IckRJRflo0M7XKQgZRXkC52ffnSczyGiMzLxBBR1Lseu
yogm0Sa9h4GMq195YwJtiNL2fwuQ+LsVfIRkdOsgMXPa5MdcUVse4DAV/AcLmKtQyRElF+WjQztcpCBlFeQLnS/9eljxCVhC6cnxPVxaVgJhWEvf0/p00iI8KGSlFlDs
/PB/EBYZgfpU0/N97hJnAj71HTn14m81fQy/PIbQNkTszal+xV0omPFBpifOS5+QCcBvhCSt5lzzPQLIGQ0EpnIHLql8/FShcQ41SVHzY3bOZQhYYNRW2V930q/5eInm
pCbms0rTz6AxWswEGdZrCtgX69cx1VQdjt/ONkfmcva+Rgtf+aIwriJGmjgpJ6RXxTeMnh6W9A0s+BtGf09Co61sSiLWde0HKUAXkMXXH86Wmhm1muT2ZIQ4GMYIL27d
YYPxyhN6SVWBQpsfvqrgkLNWftEOleNSJDN9Mtl3UivOK/7uICZb+6YHr4AEA76ND5BP6mCrLw5Z4FlvjUXCXvBqm5kOIWMPunDExAhV6n7NgysaBYBJZrSuEsAoNIeP
mdmxMTha3nvd5mR4watORuQJPeNegJnJ8HrXu1CtTys7GR+uruP1OYiIcblgqoYjbRgnWtrGwSDDMyZKnuW2U0OjDKNnsPC+k2PLs1zOjEplZCeygbXjnSw+hy7zBH0U
s9i+okYXixpSFGxvNarZ5mHapgPhbof0Ul79reLGcUVHJ8Tq29y+m4SjkExkTaoBi8PcD3kr+a9XD29sOD7MP9imIvPkNkuJfB6Z/01HJjISWdRDd6lSCnhmuyh/0wCl
XhofsD6KfO12y4mGaWLs0twvOV8SQdzWYcBa8qh4HmIjPlTJc+aE7PSzruqztFxmPzWfZUgBth+ts89Y7/+zFl4aH7A+inztdsuJhmli7NJpYKmI3vOcIRkeCIffT2Qq
2aC89lv5KWbclb/bxZxDcVWF4AOh22QSpuOWXxOft3iaOt9HGqwd3PAHZywBOrXg2uNUnV2BPE8JVrTCSlLsFYK3iE2hvWzkuaNdKXmqoltkk48UkuWZxIMQAObzVamX
oShtv3aEN2sICNFMxkP/eddbuRZNughdNWIBVKmHN3ZRutcmECTe5uvlqDEj60pzpkfjcIXcekmcXP5elyDTDCybtHT36STXU17WUSh3wjLS+vEQP9OdNhOentwSPToO
0VaekShDIf9vZWMkb7wv1ihjCialeFGfuGCGETt6jASs7+8fYucipS7edLQqcsYkuGMMYVmYPw38oSKjtJX7tIRwugVV5qoH09dInWio5zvTsO6Mk794j7Vr9iQAyHgL
3T6aBW6YuInn6neJAfx3ZzKp1zMp1Dm9NpgGMprvFNsP1j0eCFCDoEzpDXOqusRze13bIxHFqaK0I+0lu5Yc98haGRWKh2jZCqIFPXBb7FbNdL3wDZf+MHKUz5HaBXio
Ez4QP+I4c46n4nK9vdrMdv2Ij5a9xfszgEzfbV7Q/fmZtig8l0BViQbAQuw3FwOr3ZHslDznmGpU67SFKch50LF5zdgJSRwOr5glcQjS9WUCxfnE0AiPyGpIn3/t7QfY
jxBPvW3F7ncIOwB27H03cPnlccLj48NhxxrElpC4bT47EoIFdy7zAQ3E4BYvQL8SpqlX6kvOujFp9xDYVHQFJZ80OV1VfF9oD05TFD9KmiMdCcthSW1nVe5P4Z7CgX0T
irvrfLG2AAxrmt3sx757PcNGJ7RPsYRZJvniErL5An9eGh+wPop87XbLiYZpYuzSzYdAI4fc4Ltc/kfzLHCrm658g328uUACq26pFhWqP4shTDQxewMhRnrS3E+W0xP/
WvevqcPjqfSCR8VKAQQNFw3GLbjRyGvHyZcRk2P8fZ4i6LzdbPWXQ9vIM5lSymVMfIc+LFYiABY4ZQF5z855mKkLV6c2ITSDXtlPE7JMIrLe9z1qrEwZ4WloQ1nK4n2A
wZ47msNGujOSIC1pleQzE11GiQL1eHDmM2nAMdrclZ7ay7IVPQ7IO2GqYloCva4pnzpz0n9L1ryxfG84fMk6zTjnMNK/oNFevlh9P0l5fHv/tYkkhXV+DADQeGCO6DKV
nzpz0n9L1ryxfG84fMk6zcU+TUl3XBjWbf1DD7ygQgIcWdHPYxB18uMkj1Emgh2F8U8vQsJH6cdbUh1YzJNQziSj0cac0LwJYi2pgUWNvLqUJ1Ia9WeBfVq7EAYcDVfA
nzpz0n9L1ryxfG84fMk6zXHwZv59/oglSMwPujBnKk5nHvQ8Z0kVhplr4fnbawSMfX9Es0IIcMeEUy4m7v+KRmF1d+3StbN3AmzTXDOcq2mZOMOn5JyLetyERCpgFWqB
fX9Es0IIcMeEUy4m7v+KRjsAnaxwRH5+pm+ZUut0xqCiB+ev5jfjn/w9ly/Qtlz0nzpz0n9L1ryxfG84fMk6zemRzEIGtiThrjR6o0AER9i29WkaglYedFgQ84ZSHqnl
nzpz0n9L1ryxfG84fMk6zUa+SY2uk/ndwbWO7w9gcxCgXZasQWUPvZMsR/cf1fCshj/1wb31O5m136YnBb0j6ZjSDpdXbyQsfbTdsJSdPFsqyjdVeKWZ7C5NaCpXSMrA
nzpz0n9L1ryxfG84fMk6zZUooTzYA8lAilxyJZhl6k4uYpGIjaUi7tf3s84xauPrnzpz0n9L1ryxfG84fMk6zQLG1cDYEr2wWAf1i3vmiacdDzvCjNT77i2NpjkAPOm8
ME7SQwuPuIwThOITaZBeoxCJLOS+HkbD+vejgUAUYcEjqFdNS+/ooGsJ25OPs02GenmoX0Q928/S5O3KiDX/GGCsvds6uNQn3VyBx4GNCIs1Uv++FnG3jqFsfrQoKyw/
RBo7sSFDJt1hVfEuqUuVIteyg/Pwc0dqjsaplOuA14o1Uv++FnG3jqFsfrQoKyw/g/CFtMzsS745Rh865mIuyqBdlqxBZQ+9kyxH9x/V8Kys3hSP8XVY0C+l/x1OBJ4O
ggxFtgvWDFGpHlGayLAfvdJT7gQdPVMClHkI1gA5JTs1Uv++FnG3jqFsfrQoKyw/xc/x9+F28NeEWhwG+7jYxW1GRFDKQqbqBO/Mq+BRLeRepNLi2SNt5StzlzrD1gdX
qnlqtaMLIAfA/sUTElisG3bZsH84QoXIUoelJaVXQQ5epNLi2SNt5StzlzrD1gdXiewn9NQ5i/1tf0UCthyMNxdzdryIUDjmPnB2blSe6/U1Uv++FnG3jqFsfrQoKyw/
3y3MTrsIX4ahh/llyEHZiOXViEHhbuAwiyU1Wo31MLs1Uv++FnG3jqFsfrQoKyw/4C9gPon/xJbKHCKcwgn8qagPeRSiiiBSLrNM6L/oJva7sjrWKGRb9ZrliMKv+jpI
32rF+nqmF0NJ9o3uw372MAdQ7ERf08dh7txZUB8zuTc1Uv++FnG3jqFsfrQoKyw/cg19lHoTsUgWEB98EZB0Zjs+FcowHIPWZY/nMBcBQ141Uv++FnG3jqFsfrQoKyw/
x0ouf1SR9TYwKuJDe1GDI36YZkr2qoKL/GiQfrEN1/32BHRl/4eFefd0mi+YQcW3qVu6MnaBCMysuW8+bF32tJCXtHUbvcnUrHQDnnoZso6oXeV87XfBrWdoBI66C8Tt
1eLC6Jvhtty7WJfRMxP+ZKj5v9RAiVNML01oI9RIth/EmBPSk0KCZ5KTVBLjAZeBNqq4MzxG1svKKbErnAGaZJZkwb/ybModsK1wu3TIjqJrvmfC0bStZKXmrVGhpYpY
n3ZgMT390VJOCcRbkozf1f9+Iwi/SPt6VedfFOTCa2Kc9iTTwjz08rYYEy3YGEs0UOFJwZAyKwEwZu7HtI6lfCLLwxMrtW9oDHpbiHkif2Y7kja+IWUbaZ9XHSg8ZJ9z
GFzk8VbmAnvRAYfUkI32O/BiNikkTqvrnI/7A/n2gXSwv6XmLGaU/dbkr6ra9uJnImIwDeLI3c1RrYUGMzoN4KE+4rbrMMqSAjvg8ENhhNFrvmfC0bStZKXmrVGhpYpY
S9GkS88rZyCC3QD7eypI5stNAprDKFZOrSrNBnXaZRtwIDm4g9WOkPA8k3gHJGhgxJgT0pNCgmeSk1QS4wGXgfgwzH92yJ1yY96Zs7RW7QRYpDg50rC3OyDvYXlAKiqw
fIc+LFYiABY4ZQF5z855mJwDjl2NiGxw+SM9xrVQgL+olGVKtK/6ceVvqkGCMmBVOHxsjzOkqOrYiFcmhkKyW8SYE9KTQoJnkpNUEuMBl4HqZ4fr0VHrgleov0ZkYcCL
TsUB2KQBKfPbS49qhqB+NBudMUpOvEviX+pDvNsbFkmUt0nv+3wc5i5ywIcdPB9rHQ87wozU++4tjaY5ADzpvPEyQAqror2nUj3rXIObAI60ouNgomzjPv4xDxjaN1sj
rGj7Bz4pv9GrDa7ZN4BnwLscyheMGBf297+1s5w5SCMv5Kv04pJH+da3Szq5HHDqUpEJcA+JoTc5gSn25PctGNCGouRUhclHR/INQWyPo86dHUaSCpbKcxFrjfw8aQ5F
T4o+ycFjNLai+e5fFZWDz15Fkq7cATSGA4TwcTPzJLXmX66+R0zaUgZSISUqUQD5m4OEJ2pcb0ehjWXgJxfpwVdE31lvlpdd+LiceupMmJzSuEU10ThtZXIMIGbqzZbZ
iY1Onv3JhWzY+O4XzF4dg6LXSKOX4ZP+zyikVPVxrce3i2idn+4+yAXWCD9twfyrPZJsdnIIKaV1ENpMvtxHS1Gi8K+QXQ+b0ucrpT9/ntPuJ2j5kfv3NEnOkSi6rl1o
KkHTYLZ3eFVgR6Fcq8b8rDAimnH+aRQlrvOYIXdnXYIClpM3ZnbYwgsUfw37V4EsiW90qW1/KeSF6cFJd/LkPokPhgQYYiJle49hR0lQuldWxn86rTgSwwaRfzq/vXfA
sM+sLOC3yGjoxPGgBo+9iRf+Mm1rViRwKJhhP7jiXyjmjYZGTPpx5fHkDH12aeTGdQ3Q/r/Jb1uhGcmKkH+fiVEJN8Jhh4pj3pLNn3sJep8qQdNgtnd4VWBHoVyrxvys
+o67C0Xe9YQdI8Z462KWH4hRfQYi3US3QdbT3igOStaD6/lRQnJzuhZslyegD3NpG321qrp1x3RvakqGaVpErN5Wn/1K+XTf9v4tVRmqPDphN3Oo+xyqSdgbFVthU1UC
ntF91Ls8yxOWxYI02xhwNHjFf+6q3fiC/j3/JD86jmqjvYC11sLSYDNzax74k1xJY9ei6ZMPDfc9kcidxtiLnFYG4PBB2JSr75ctCGehM857zPWXQVbvOXb0cng2PVfT
knPuxZJ+NhY2VkIka/CHPJNQjfB/yCV/QSygCHGXPQgGbEGvHl4i/X5gaayJ6Tnve8z1l0FW7zl29HJ4Nj1X02Jg+GqCgAI93a/1uMKnMnyUMWO0dpQXlkFdMtf4W0MC
0aJzirHh5e5WbaruMV0duSoXIDoGUGpKrnKpfHmWyX0IbwKhTJdkXICM7eD2yr1cjANhtQxAL1JouMqBLsG6nfUkiaaOwGYmh2dHj1iFzDCRYjIQEh9DisJEJ/SSVF7/
lHBEs381QoTzd3jX0UKdfFCVWohiblEguugfXZpcKH70U58uX29e53lbBwx48mpERVv5Z5X6Ilk/J/AtTlFDuKVwtUTZJC08KN/LgrfQXxKbU3zzgo6BuFtHJe9mwMcn
Gf1zPlbMWClRNWPsQXI1F9Q7I1CFZs41TiJHnzmj2/iGFXEUKqWA8GGrEsIdBR0vo2EIcBbUVTUvp8NnXtwPDEIfXJCV8KDZM40hbdm02TSP0lz2vnnCJ0Tn/Tz1lTsn
FGxIHO03SLeFveR7yYigcGs/2YdnU/+gXkfvDVvRqQK4xGser5bAPhNbMi8xmh/yhjA5LiDgr++DW4qNcM+tPA2gDC91L7Yl00ArQmKhMKcytN05TBWeeR1FG8YqISTh
nzpz0n9L1ryxfG84fMk6zWjNpsHcowlWOTEBVCeXn2FxLod1BiSWHo5Za/cR8xlTH7qsns+3drobOr+zOqQIW0PXMd6b81Qq4WmpPD6JFrY+3562Qfdq46CGPZbry5PX
UNsLpdcB/Rq+FRHEN6BfqjlD8PE4aTVxlwqqgna1Uqn9PcAmGzWops2py73qK9iNn2TPuABIPv2vzp8UBXRFQe/dGDcAx6P0tSH3SjheRY7GCZHN/fAWYl7JJRsWJO01
B5tDItU87VDrtayRjNN6dYrfHtgFEAbnlv6mia5w8W0fuqyez7d2uhs6v7M6pAhbTBqea00X8Xh6DcL7E3P2sOA0DGJAbPFvcSuKDjDji1Vf0quD23WiuWLKw4HLqRUv
a09mi2KxPKPeDPEacp/TAI0iKqWWXEKTpEiOJx1380lVMRX6uXEvY1GGvxg4T4RqaCTcDN4+BsN8FnupQOVKJB0DSOseO+pj5mYM2GixL1uyK+DZwTG60hQlcXbhuqNB
4yPtqC0rXF92obofMM6Zue8voHdWoEV7zHhMeU3UohmdLNGs4+HiCIOWJbr6dfVbPt+etkH3auOghj2W68uT1yHHtdB3nGDPBcKy0vTvAte3Zh+cW4mI18FQ4H0Ie16L
xGOGMOu8BoazpBtDkChvwqFLeDrG5p3Yqv96avuktoAytN05TBWeeR1FG8YqISThnzpz0n9L1ryxfG84fMk6zWEU3Tg/75k5y6nVpcAiPfJJQtdiRpJbCh1Ax37hrxbL
H7qsns+3drobOr+zOqQIWwimVm4kqQg+Ty3kVjWkWPRhJCiU/uxEu9UDk4UIFrYEwkByTZojkziKZXoORqK6aQ4EVXxMO+wrOkxR65uIbZKh6OcizF+Aj1ZZFs8AeCnc
wMjESQuiynqNTmFhgubNugzHywa80PrPdsVl+TBS7vAvcNOislCAvv2wC0lpnAScaf/qbUXyexoOKDf3YN6xgEFINYaRRTXWMpOA5GwHqBofuqyez7d2uhs6v7M6pAhb
jFtykjkmGGpRFy7vOCtYF4NpYs+SMViUyyWDxXrzCZraQNj/5kB0kx/RJDK+U+ZFrN4Uj/F1WNAvpf8dTgSeDn2bStwbsT/G5CZc+OiwMdQJYdgqs/1XlJDHD0r867dY
qpYTK5hNmd2Klzfb/6YEmYY/9cG99TuZtd+mJwW9I+lDZfZjH9SyxJ9BrWomFmd/DCPNmB3/RMuUbrfzOZJ1DoAOnYg8ewLwIe5dANcZXCUwotkTZHj/HqDH6k15j3s+
LpsPj5eVa9rqn6CY/HuQCIhfT3O3II0NufX5ovZ0IrfSx8btrguOvnXUododCCoFxOuLF8bFCdc6wlwVqk2A626HBwSEBz6S1h7xEzoqQSinphJRwnK06j6eR0SBJ2uM
g3nLNqYecga8utXofv3f0cqFwZtCdaoT031VQm6NB+0EgvAM2/L0inFNwBGDtBpgngju5HfLuUTeJAcmmqF0xt6qxE49samevIi8TBwKMWs4vhthuYayWiToxMRIcMJk
9hro0hnXZa4uiA2Smr7fMDKGVpAS5u4SzPYEcIWxB8PDnzXbEnhyM7GIeSfXUqyYqL8yhZjeNPODdF5jTxxiNPD1B68uB8LQA/kuQ+NtD7r0TuTIdP4pGfs8VHXvbq/l
sO4NKE5LmIKWwaudBjBBVXl6yzhVLlcXtxiohkB0h/MfbN59wY8VOUoavAEO+k4AF+WORhXAa8tUnw6+BXnVpZqV1L1tNMrd/sdf3rOrhV3lM60Oai5rPqgvex2naxP/
QgSb1hr5OwlNXbJSZ2/PoiBLJ0HgHIQ9QLFOEoxkbarbQaiylWIywYHB7ynyk+kCjPkZ9VafcuTlwxme+WqeMLDMQkKJbuyQYFTmsE+qz5TIBqgOraBMgPc5pH1OvH8F
Ym7g4njev+mCxidod3fMkjksXErSLqd0lQoAzuVq3Hsnu8ZBYr3GwwiJDls8bZWOkI7xdMtKa9tRu/KT/MrX9TLyL5SjU32GDAOtHRVSCXB8+aDV46yslnzQlZ6CG4nz
ayCV4X8QTuxONsfkr/eTslzvXxZ+J2NvyD4xzVS8Iuqqiq3WEdnEpA52Lhw5PbJTn7zO9RWwNrVt6NEBWsNIAeY9wofYoU0er6HUrtwhnRrUgcyDVvDwzjtIkqkGkLWp
2UVqiAOBE9mij7HbjnWR9Pz5bGLbzOvxQG/tdbv0FC0dDzvCjNT77i2NpjkAPOm8rcA/X4vme09lIr6AbG1JZw/9166IQOkd42L7EISGfva0ah3bjQWDS6/45tzlep7D
rcA/X4vme09lIr6AbG1JZ7kFNNw0xEq+4jre/PG9io8dDzvCjNT77i2NpjkAPOm8rcA/X4vme09lIr6AbG1JZ2RROeZfSM6kcsLR0Bw1JfS0ah3bjQWDS6/45tzlep7D
rcA/X4vme09lIr6AbG1JZzLyVTR/y+LPVc5yLtV550S8eMDU3kwq8F6AsCz++QZzL1xpWNQRXXX6GNUOqTrtu8ZD2vVscriFeMhYwB+ZTqpkjb7owkbC60XvVJHOWzyU
RYW48Ty988nDAMT7wBLmBG6sMR2Msv/Iogh8c636r87ZFJEYVKbtccWGJl2WYCTtzKHK/fHQkyrtMcwwRT64Dz8QOK4ej3NXDlHuZTnQJao7PhXKMByD1mWP5zAXAUNe
AdYwkQhi0ByswG87w1GPBjaFBlQDvL3LJjFMzBgrR5R+mGZK9qqCi/xokH6xDdf9zKHK/fHQkyrtMcwwRT64D8WN41AojTHZrhrK0EVAmi9grL3bOrjUJ91cgceBjQiL
AdYwkQhi0ByswG87w1GPBhPaPyV+WBl3H5vL3sN6D5+VJdnyU/Dre8ETDdm/hv+brwzArZSsp1dllT5X56n2bHRFID6U8eWcaAm6cPKvO8qWZMG/8mzKHbCtcLt0yI6i
rxM4T7cc4yoRD1G3pb2xjXHzghdMIbJedTNKiWQq/xkIAooEu/JTNocuNZb+KA5BFR8GFkJo1LBTThPEHxeRISDQq2tCAni2FqmAvCkRnd6upA8gxkdCp4jUkK51DgVi
m5Nwg1PyP86Tk/x1eb9taLBtHGu1IQjt4yop0XPVJvq0ah3bjQWDS6/45tzlep7DeFcvM1hgJtWOCufUyE5B22ROSutvVZfbYnzaDS7IEA35LC1RbL4NY0NsTaUbf6a2
Oz4VyjAcg9Zlj+cwFwFDXgHWMJEIYtAcrMBvO8NRjwbnUzF0bz0GUkNnQSEroOB7mHvRt3HwAGy2sgPH7A3SkS5ikYiNpSLu1/ezzjFq4+uGxQKaqYbl5JKD/vw/je77
XNl2sgqdCMBE1ajEHVYIxUyxa/YnDzC50glAexdmmo/J6cS9cy1GI4KS5HU68ZdwcfOCF0whsl51M0qJZCr/GbDzhv3gUKasSx3IKjjGkxWb2BNh55TQk+b8gwIF7NFp
MNbAH5bC+b+CLeuO6OaUJjZIpe19L0WIUbxsC3TkDeYLjIYLOQwsgvz4rXyFXgV/DaCxRn5y2rEHEv9pMyZqixvkgnqBhpdTa+5nfUO85oadJR9t2dXzCIrOJ+IqzUw7
1I0Nog1MHkzczHLlcSNNWNkUkRhUpu1xxYYmXZZgJO3Mocr98dCTKu0xzDBFPrgPG8RefSLl7gXP+rof5FMJFkrO29uyIkswek0FoLPfcUUdDzvCjNT77i2NpjkAPOm8
hsUCmqmG5eSSg/78P43u+2912bCXYvnMs5EaUus66YxrjkBAT4K9Fu0Qt/XM+emirwzArZSsp1dllT5X56n2bNL6MDDIKyL30KeBU7AUFTxkjb7owkbC60XvVJHOWzyU
lCNmu1KZT3Tk2cotNgOUz0ufTxSsvqF0/FCzYiM3SCx0m4EEG9mVJ17dWE5OAOZ/Zz91t8pSnF2TK/cVa5jTfShvyMm0YRf0lPFb5YmAziOb2BNh55TQk+b8gwIF7NFp
MNbAH5bC+b+CLeuO6OaUJjqZkZukrLgaIFKZrbGIuQT6bFDAYBF/dA7tw5u9g+oShPijzFSxI34OyKKhYOmhXQP7mkwPIC9yuXtVFQM3R9K+JG6zzXZift5o3lAtSV8x
BfHKrlqMjn2lCcHNCbhNGEWXe12JNl80i5wU1R388IhB58nPzQkRw9xA/iA8ZTYpozHrxhHbHTlBDg3H+hrn1ap1sygJUJQ3Tv+H0WLNLEWKN2VpvMrgxGAg3TTfmvsF
rxM4T7cc4yoRD1G3pb2xjcJzpcM0gUzoVEjNmX6mT1NuiqyZR4c20sSPg9f0Nn3eYM19dYvShFdh13e+CmA7OcxapJACFCePTXgO73znTh8avfgJAtYECvxHOE0aRcY+
b2c/FhwgFm76cayrLhJAP5QjZrtSmU905NnKLTYDlM/zOZoNt620X19A0E4aVMbCJ1K3N1j6QgMIT1QUZReHe2sKDbt6FRyZTA7OrPDLSbM1191b0jbD9Vi90/0jHXWq
nRYHJoaFQXpzmHjVSzUVSKanmPgGDdGwgaUf8jabfg3lb6rVLD5Ox6IjmPgOoV7vWAX0aSq8jdPnfYofg3WoHYT4o8xUsSN+DsiioWDpoV0hsjjUWIWmKYPITa/lbY2T
IdzUELr6OGN8CA5vDjFYUcUIBeuk+1e2JXKyMF9BpXPWr0tBa+bN/X1oQ3I8FThmCiwHhy3ClQmFIDmNbu+0klEQu/qP4fpGHrE7O/IqAeib2BNh55TQk+b8gwIF7NFp
2+iJra9EvgHQ05JXSvuRIngVRt0RGzFVQGKmeAE4aoJ3S+ifYHNyo3eYkwXhbqYpCuWSSEZDp3Q/xaaLaKMb2QhIdVE/1j/WSIM4j90pbJ4JAzq+icl7D/wDHBcj67+8
FR8GFkJo1LBTThPEHxeRIUjyO6wFpfx6kbNsb93UVmvusK1ZMYTi5AugxdSAIQWzy00CmsMoVk6tKs0GddplG04lGJs9AtxpJkcCbH2k/Nu4BJXQ70QUa0+puF/S4lgl
EDPck4cqX5IMI+p0nK90op9iU7dSvKNRmkMSXC0tbOh33Q8G/cQi467J2wCaIN5VG1PIT24vLdYrqg/F8N+EHXSbgQQb2ZUnXt1YTk4A5n/mNcKjyVvA4RBSrp9kS42I
k03fc6PYF2nNoppX1YZC/Sf7LGykourMo9yfPPGXIvAsTyMnDhNFLppk8CSAbu0X2RSRGFSm7XHFhiZdlmAk7VDfG+pWVic/ETEpL1c2A65QsIRnbq+86r59p1VtwlNM
0a/m65fad5LOU7q5oQGA3UfrE7FK5jHQMBNp2BETaLaw6HB5KqAOlgAUNYUkzPNbu+ZvXVVv1m5M8vs1fbL1HdjZY0ooxheVQ1i6IMEEfEFeRZKu3AE0hgOE8HEz8yS1
6kMkZ3Lq5ERp2HPxPzbxrMLzxR6tRTGMYww6a1evAzGpqdZqCzNN7n4cqeOsizSrKkHTYLZ3eFVgR6Fcq8b8rKm6zDCoHBIi66y1BSXPSrrCeGlVO/DCgmv9+0YTEOIT
ZOxoRqZYLELS36eM51O3yePYpK9igx5sBhjqKI3uvc+HPjir6VdAi1Vd2Vy1GdA3R9pYgP+eUaTyniPa9xpysDFiZ/1N++J5mriLX7iVoF4XaxjxWybuGefm00d0qcKy
T4o+ycFjNLai+e5fFZWDz/rTwf3ewIT8hWElR01ZUAUIzY8WUmwy5FiGK9hPwvI4ZupDIWHg8qsDBhhhqkznQGzSgG42esB4IGN6x9320k7s8zpxvNX1mlF9vvZuZMb3
HDYagQiBZ4EehbTcUAYSvenm5i+2h/PiNvu3x3SUTuKT7cXh608zlLg+N6we77EO49ikr2KDHmwGGOooje69z+2w1SP1KgiEm6NTzdyQ5raPZ42TjVIRYyJJ5wVspFM5
rZY+XdSkH4lY6omSSWNTV6+RPaAi0JZS2eIk/L+X31bKiCbRJr2HgYyrX3ljAm2IQCVCIl1VzrT2DvPr/xIXDMHQUw/7OizKTIILRdYtbbjRFqaiXdT5BU/1mCEp7qY6
jG1ICoUXifFzWooSvonvwsqIJtEmvYeBjKtfeWMCbYgsmE76KvCsg6TShn1bmD6GukY+Nab1N3bXGt3hJOx+Wll14Z4lTIZO3gHYfBLAY1PArbjOPNLQA/v2SG3tZ+xx
e4u2tEAk7uRQBfIdIDgMkRM49mSZXXN5cvgKyZ7MrzL3mg8iw8phEXkMSay9z4j6JV5BKL075q/MHFGFLG+SHmtr4vTdN20XoOZejtkfvzEPWjHI+UtybbSn9Xay81MN
abTNsrnFNtuHqpYL+jQ180TVHUxc+rRQru0DtZW/f1Ymbm09EBz8e9Ix0hWeEvaeXu5JF0Jk/bHvHirEkP6tnRW67WDOVl4ibXuzXIj49D+OFbs+ZqprkBUMciOgQlHV
FsF25LkAhyxrZDUUBAO0pCDXG3omaCaA0nwKOxpAaE59pQar/H2x2rixj+ZLfh6CwPtLJ2oEHFBGI0Y1vK8XkDqXqJNSNfqgc1JJEpnygiwapCyFy131BhHi9uUtOlxD
ghVVLdbo6yNQLlrBboz4TZiSXr6ucnn+z4GFgk4ov3e+BU+n2kb1+U1pv9l/cUyyita9gj5lX3+ve1KzYXAoPRv9EtMKxKvJG1loG+gEuS1E1R1MXPq0UK7tA7WVv39W
zVBZPCYUjFwMnZXtmmlcs41OmxxR1floY+PsihJkwNZXDH4OzChLhvbqmLXvhM1DuZ7TEdmSZh+u5kJ6IzVB0vT1FusBDHrMHRO9wf4ahIbMcBl94du37J2x4g6ki+k4
msmERYoybiOsutPrbhjvPdreLSrfxTLmvUjdO8YCkj+Rzt1dgNpD7igdalnx3m/8gDFgqQZLxM/qB4Kt34+db+RsiX9boD4zIfwpZtAJ1ZqEdWC1oKIGUNDRWE7Pm+jo
LeLKo+D/s4lFQ3t/SrnV7dEQ4ZLkDAHZGl+qouvHXfDEvCElc3Vm1Ppw7MUPzsruYVyWSJVi7CbOYFHjrAjUwE08niQdv22vn73az4dpcZx/3re3cTkfgp46/VJ36Ozy
eO+d2NVvnsHb+1aZ6G9rqzQh96RpHwsYhxtCQDt0FceKrHOo8k4juYCZzzL/vTX7QsvRoPH9poDPRCHZV3pZWVh4Bvsxvhoizsl6XT0mWWujA4flyOWLfuEDU51h/ly9
eO+d2NVvnsHb+1aZ6G9rq8CZu6ZR//0Si5dx8ho5miynr2LuqM+SIzvB3zE7xv7eSjPA2YAb/WyYcBc7C0jjHmCVIDN6HyZKcSszOefMJKTe2DfolkiNM3wPtVD1H9Wy
2j3pAtgYpKfwypUScekngQ330KI0dDz2I2FeuGmgqcdI0oIBOgZv63DdEx+dDnfW7clLDiQ9wkvOWu0syLAhOyIvjb/HX3gDbhrHdYmkkmdhgxuMmCAs9C1896MHOOsa
RxXvXL7DUygGwavjb/FSiG/ZLjZLyFovjCB5xkR7rZwuOAzAnb+ELwviN9bPoahBpSt8RTyfB3WuXNq3V4YX6EHv7wuZNvgGQDBLgloty1dHbE8R0jHvFGkRAPbPyPGB
WuEiOdHZkRf3lW1reBJnzPCGPNhqLcADh+qUVl+Qu3HLwP4MkH/gStukYRFN+q+XD3n325gmAMc3/imIJPP3aqxo+wc+Kb/Rqw2u2TeAZ8AnPUyPFVX8cKpO+ySb+a3I
5uvXTHafDiFCwy4B8p35N0+KPsnBYzS2ovnuXxWVg8/D87qY/PprlKgpuEs8lIACbnmxuzIELf2kQi7LLa5NLSZnib9W66tg7Svh09ur86KUuU9onqco1JUkN2DVaGmu
iDykPge2eUW3RxMBbR8zBh7jD8NWkvjFWceQgzOhgAF/WM/VJQ5ep1nWYtshQ1yIfVrzc0ZZ34+1QRt/XPvngfCp4ipRK/eyh1TuJ5Z434E5QwC/KmSU1wJkC4A/4bKG
RuRBWfaEbNKnMHOARDgjNsJ4aVU78MKCa/37RhMQ4hMucZgnqYPZnAO00Dss/gtcxnkZHuZblQ7kWJN8UbCuYLVwuNSAvrQ7fUAyN5x1L4LvcBV3RMC86pZ//apWOIqs
4bg52vsr88MsxfKNXfkMdUn8DVntKKFO1smmDfJUjtySdV8WKSeAgcySCyC4TB7H2LgyA+gBJR8J2jNyxFdmFsYZhaf2XIzJitEc6aEgvZKKvtUVRneGXFgUF4MmESWi
jOWabKrLaEgOwy3E/mYi8ifZcsbr8AS0IXcujMUDRif4PwUsnv5S7EfQqCRfx5rPdrfKCSbPiRbydA1yTFKQxT8TOuyONEAISEY1Cy+mmdHUVEU/ZbschZglUkmLxhBZ
UaLwr5BdD5vS5yulP3+e01hMfxgkPOTdyDjVGuNEZJKTXVKFNFNisvvk+illDBR1zfoMmP8iZ2JkvqqilftGrBe8OITqu+QLvSbN+ApNFDpzBwTsakwsbJW67wJ41pxT
yogm0Sa9h4GMq195YwJtiAx1gG5LuxSVx6d93HZEIfIUYCGzV5x5Du0hAp8oNVhEZJuKd4gs9a9GXF4QGBsKNlybRzfqYMaJOHPmy0OQAS/VyHaaxuY//radYPPZjdTb
ir7VFUZ3hlxYFBeDJhElogbiONG1cvLRggNRnkjFIPAoZ1kk5hcmwXP8POW7Wg4ryP4xsJDQN5QCUzHwO/v/Kyctb/lNfToPmYAhOk6kc1A2AFpkqbBABxAx8xEaprRe
yP4xsJDQN5QCUzHwO/v/K/PZv/8pChv41qYO+IfBNRA5a39oVwlTdcxCW7tiDXVMUF6AGWIK2T9zx5IbYcbM5yGttWbL8KLF4TyeBF4m7briHj0rTxoZ6bRub8ATr+vm
0VE01QtlmbqxD/YCqibXe9TQ6uBIzLMUFqNP3KJ722fiHj0rTxoZ6bRub8ATr+vm0VE01QtlmbqxD/YCqibXe9FEloCu53f0K5WjeFpQSBcVuu1gzlZeIm17s1yI+PQ/
0VE01QtlmbqxD/YCqibXez8DDYlKSj6C/ZHIzniAXNhxakMIeJ+UraRTIcOD7H7AJUxFjxLT0tV5qGavxxn68qF5pTS00U6goRHubdETP/HBrwZZAbTiws17NmKj98u+
jc865/9khik+u7ZjLhCnSBdZz7XO2kpNOdZWIqQfHIS66m6GqTyl3QyMJrfh4YB/2bvyni6QJfRdlGFoMI7h8txAtAPzpDMZ7ktzKzGMALaTKM1u+2Wg4xOxaWGRQL5K
bhft4JEdJ0mV7Trz70SUjuFEhPr4QDHD72JTOFMc++EUn89S+Y8Lc/Od9iO0B9vDhB93Ve0L3ybxlDQ76FnDLKGu6nvMYSL7QJIqSfEO0dqns8NHdjat5DL8rUIdRX7/
ZJuKd4gs9a9GXF4QGBsKNqHcCDYOhXS3td9lFrGLylg5a39oVwlTdcxCW7tiDXVM5jOhgiYF2eYyJas0btQV24Y61d4LPPRH+yWQ/igCZrbKiCbRJr2HgYyrX3ljAm2I
gscDtCgzeUlrYYmBOD0XVvY1Wxtb/+HCU8sayRAkTbQ7tHiljXORXyEbcRzJwL67bmcv6d0/zaB7yjXwbh9Bh1fcnZIqyB2M6Jhw5Egm4joyy664+N6Vtq2lENsl/h4I
CI1tOId2H5n1rPKsPI4MeN3bpdWPPdpQ9FzpLQ3HVzi0Y9TPo9zhkIiXwTe4GYxq0kxnjm7O3yvR/8xOiJwUOUX2YPAgRCEXmVqyWKzkOTbIQ8fsjkVZ/YxVzddR7bnR
RCKdIPDiaW3782lgue6/NeZfrr5HTNpSBlIhJSpRAPm3uxC1G/9rDclBDv6hd8xwEfSqTYzX7GjfVksxwSsVjsqIJtEmvYeBjKtfeWMCbYgn3Ndf7YN1AueBSy607aa4
KUp4Ohv/R//n2/QtfcE/Cs1NN34imNs/Zw485pjQKsyplHO/oimgxfmeiuRceW1qLc79V/vlmWO6ofuCX4ouH0gt0CuBCVypwWsnm0QaA4YQPbs9cKRIA7SzepFqQ+ju
KkHTYLZ3eFVgR6Fcq8b8rJgcI7XgxjbUQDjjb4z1hVXJatMs5YEpHGpo7spmx2O8m5WAoMyO0FfVU7zMGB2kGshDx+yORVn9jFXN11HtudG3V3odZvGMXvx0QfsQBGB6
cUeDM9j+eN5xMsB0EXmiwEtNhQS4UzOUU3TqVu/vi3enUJs7QSurkVb5vroxCe3vHTkqAc4Juof862wgk9NHO8b7ofViAPZiqc6pC9jeG5t7AT7xcfCrW64S6WFL13rq
AIrUifyMVWfBVBKCyzJDMqiTITm3DKM0xWs6eZ4BIf02xpM7WdSBltGnXBOj2gfkDkNlpL/ORqZzJC86+f+l9kJTrHBjyPo3ItC0tMvr9p1S1zAnlZma5TUNAOnhrX3N
cmQrjzFw1u7gEjq1kQ4xiDbGkztZ1IGW0adcE6PaB+TyojDWn8TkyIiDzHndTx/sQlOscGPI+jci0LS0y+v2nTUlPbu/IJODN0fSTENA+llR1VmSKxYVk+mOeS41IchN
lk2yctemLPQj8x/MMiCtpgMWO6NgcgDUUln+5uhF9KVjuMmzOUM0aZYfLq+BC+g9LDTuwOZv2rY8j4iPikBrfwaVXIy4NbhrH3Qi+t9/NGLJl9PdFsLnVEyKvFpaRL/t
g8OhT5svMVDdv5w9gKLYlGEGnnkYsW0FlxIfRrHbscq9tCS8hc10KuGHhiu16GXrFec2qryryekze9aspkUEmW16/seXuT2IMLXgt9d60SpD9crDsk12/xY/QW6YIjVp
EJbN/yA36kH7SCjXFVpYd7Nlm7CJbJsmq9avAIiZ1omS14yTwdBRGUf14Lz3XOFU5KxaBa1lKiut1DgD//LhafM5mg23rbRfX0DQThpUxsJqYOBtcIigFosr4x/toG9W
d6Njs4ALQnWPUVT4wU6J6bMdPnzWQ9dXFVPkE00W6oMQuOjZCdCGQaxFdPV7djS5CdTQc2ynWV9XeuaD7axxwFf3zHFPUq0ZbuWRihQMeAjnNo5araXzMixfGRn4dS6r
KnwRiUY8HBAkkKHjNnjtrSMxlr3fI7eTX3H2wbR3fLU/2ZkdW7aiVwQacKfEBpWz9D+wFUMQGJHWFtZ/fwMiMyhFq38xa6eKEOdzG+FGY7kBkpdh+ldxG6KgTxr4iz/F
Z0oDFLS2SG+SkJ2nsnjRFuCuLqYyol01G7UVA3l2YgFkNy7L3mku0tP8VJd4FfmQq/1U9g4D/tfKFn2lYld8lSX5WVQ+KfyLeHo+bY/tBtiB8WG1Rf59oMh+hCgYXgVo
UyVtj/HK5Nacy0zoJ8qsouLTh81TdYvpNLiSi9f/zTiIGeX0A9Y4DUur+JdxQ9ARSv7rAU45H75SxglG/qHxhcNxh6iYjLeMFiagP1YkASk+khxEMw9VmqZRTU4FgjN6
rW+JYTcb9fa00VsfNbKv4AGe2hw2iWHe9qkZYC0HQK4WwXbkuQCHLGtkNRQEA7SkYTGsa/bMpOKRu+06dKtPtu8azzcZ+vlhTef8H/riY7eSiq6nrH0QV6sR0TyFsX3d
7xrPNxn6+WFN5/wf+uJjt+y5noi2GjhM38KS5COqFqyNcwT5ExRmJ0o2CM9dMmtQjMGRJzlB5bTr3zm7lFOiqj4mcjL/cnBVtDxLfXknxBYCZ0rsP71dWysVQ2blC7zS
dpsWrei6oMGhXuJdEXvTmhz3/GQoGvPYzWsQ+rML53vTYCWwVj5yDVdtizfGb1VdcDtYW21g1URLnkAyJ8MU2fCrvgai456Dxs1QJVQjcviKq4jLhNg8JCKqr+RqUeYU
zTVD5mLc7fZKi8lTsBoWeGkvCu7oYHlcao6NUisG2y8I8kRLm3e8Ab29BuZOlCVL8NdrBGxhbglQPwSlMRPAk17c9nxWnMVCweRXox7A/iFycPFY9ogtOHx8z/sVKJvp
GrnATvVsHgXvHMrFWeReyjnBYaI1pIYDpKly5k2U7/rbX7cEQLmDyjjf8BuxlQx1Ah/N78V/0Fjav/9nKzdIp7Sk8BoRgDJ04Yv60TG1cr3FvJxrhCtNsiImEMLgIX6d
hUtOs3aIVSwTxTJtzRnvn+COTlWICdTDuk5EuMnFRhDzFK7UrcQOCE2lOihTC4ZYV20iCs/NRu0sYKPw8ahhpJwZBeVv4ZuNCmR23Sd4W8kSFMByRr9lVsYdbyRLzdrS
/zOQxAKGvzZStvXO4qv3It01eFtNVhj1KzSUFz+kf3gSso1WMQ/aHIaOWg7LfzkJbjFtsS9isp2PK9xEbf3Wed52Dq92wc+T9XHd/8JAytBWBX4vFGcEwJ3QFdOUhb8I
9WnUPe6zopxbEa9XhzaPWadM5lMxOstOJATmE7zdnVYEBUaI9JMA1mSb5IP59QFm89p88/lw7yjgUWBPJY6IwEPbqN0QDnow+8j5BayNcGW15V+rLxdw2LEBBDdYIDIp
w5812xJ4cjOxiHkn11KsmPLpGGvhhp9driM2ZrPh2dRyKYJBLltwf30IZsadUjOygamJvyarC64CiovuaAyh6LCgVyvCtnc0UOYn/XS9JumtsUY/X5/8+dAmQeErpkUz
vL8C+K1X1lb7aYX+p1r4Xl8sz+uIApomi8Ukr0tpSmIPWjHI+UtybbSn9Xay81MNT3NwB5QhbFA8AqzJ/4aKrsS7/4xbO907XopFvGCdjtqDEsZ8KRCveGtl82CfFsvV
sHfRLDM2I3DmS3xRFnkixPyAN1gAuN569dHrGsLDydk2xpM7WdSBltGnXBOj2gfkB0nRME8mfi4PvgX9pqzDVftLVcciHvbp3STllaPeNrkT4qNYwCF+qcROxIlqxr/J
FwT6p5yZ5zk2x3A04QV1ZC6n2vvXOXBNPWPV+1sIckn9N6M715HulCLBmYhgdZTu8vHJNmqGXEHnutvjvbOhHbp+t60UbXvWtEN03/g+hQvNUCeYVNI+4AcYlvX/R1vF
4amgdiW0TbgTHURJLxddWPLpGGvhhp9driM2ZrPh2dRWvDfJBvAl21YbzbPV3XpjI1M4XhgC/Lh60PhOHlRdD3FkvBgylHjMjP3dDsJgWJynALXRo3MiBnfcYzpwWnlM
XsAgJshaYFLODtBvG/hm7Y0F6VyqRGjw3XkOF5qRjoJODivNs0cHRLiZbvFGR75WOfgK+fqHAQ07qyk7qNJ3XiRx/BBkgvZNDlehtXNmVM/Tr1miqgs+nP3luj8dkeju
WGQQEZi2V3pLD7oBUbsE0MYUTR94u03TdurGdPmuBMWHXvCmyCNhGa9OEvoO3FSlvCq1OWrvJGBRAT+RjfdjdTbPlWEY9LyY5vK3BOKIBQcX8nqoCLTIF+RIwdrGwWGD
lVZ1JL76nn4PPd3m3rgu8Lz7IxHgM1TgOJD8xQgEcjIjUzheGAL8uHrQ+E4eVF0Pjz9Y+Ci27W2u1xVFi4wRDNynGNtO0SyBEE/lnZbnnwL6TKnsRDdUgZETqEJiDdrM
laVSsdyJi16WXcKZbNgid2WmCSUcT2wfbnUY8/+kMG+UqQ09bpKC51tpVLEj/ri0LeAvh4CT3gKsLfgs6MCJkfsv/i4O+Z5MDVYuRQwXWmv0EcGyU5KAZBYfeFSZKHlo
pQBnNmd1rCjcnhdWcHMdI7TXKDoeHZM4JbTtoIJaAyjR9vf7rICwMQjq5hsCq3IdORgU6KN+GOHYaH3eY9MhDT7dmFQ5N4LXEf2rkwKgcEswl9WAWtwaMis/03Sqez4h
OYnZ/JpcK0tlbpiswdw7+6wjTeEQzO+Izw+haGiNXaGOUWZM8tb/xit/2hbdLM9J62ZqZaOzmegBPf62Gly6Mogv1EQyK/1tNMC88dZrUtwteeE73sZvFDjytAYPsNqw
T6dseWMRCNFVF79gqkC/8wzCRUY42K859XISdfvfWK2QuUQ0dQFNg1Q5JkFUKnGHrpUca5jTDHb2iGh09ckNKeoQrQbkZ5GrwxcjGxNosygEzc8gNNjz1kx9ObQdGBcv
d7LXpa5M4tNcOnZEK2/rGI3i5SF7FzV+TmqyxXlVkkp2UaZojsTt0P2QRjlQc8qwuBfboL0qU8999Bbfpgi8iUnWNCDbsM9F1RR1t1T6vkEDp4FKRX2R4nnf3nYY1+rp
SvhgD/5uSLIqHZLLSkyI0nJw8Vj2iC04fHzP+xUom+lWSnO4Kix7StHPFd9qo5yJYEDU3H8z7GWcNAsJ2iQ8kt9R2pkt42ma8k5YO0r0bz75zDxQYXYfkeUcdjWneTRC
pfp4QYd1vAj9Wy5rk0NbrbF4HVpgESGnMVkF41EsMcmOC88ABZf9UzRlnaUbdHUXm4ZOMhfVMHthB6UgbjtapoXnrF92RFGhH1klDGRNafYluDIxdxX0xfgHrhzSngxQ
25J4qVed6UhW4sESRbIvYlSJE/vWjhz7inmRLDDC5SPFFFnXnj558hntajl6Dhiaygp0kpwlfmBnswhhLkXkZH1A99xj0r8yiY4kWvALi/iRiW7+Eo6wT1rY5avks8Li
AhdvcryAH1acFVsxirHChPInP5mL+sZyAXyzVFo+qbkd/UbySCKYE2qxzhD76n+YKKDL9W8h/qWxTQJnRRrV1erB7FwyGnFeaQ6w8sHwuqj6TKnsRDdUgZETqEJiDdrM
laVSsdyJi16WXcKZbNgid8JoUjqx0RYb8boAoJKRVGUvVHEkvHdqdCNQ3VFAtr51DM7x56GHPDSe9AzHDsU/PPgqMlGFJlov4/rgt21PvCBk4v9qt6V9k0Of6u2r7jsj
CeqkT+wEnHaMVat2nguc3ouFVsLhXHYr7ifXRiMqw+SrLlVeQDqb2DrnzVo68Tq7qmYH9Uq7tL4DLSSHqhKTG/Icu+TcSt6QbREAaBK3c4a+knqwiN05f8vamm7JebPn
uKq0GQ3MFrow3LsEfhVKFd0kTaTCQBy08/zBI9TnYWBsC/L/c3ht0sddO0N2y0MRjhW7Pmaqa5AVDHIjoEJR1TLzxmOlIy5O+FdmAVjG8KWv3CGVZMrzlxbSnDeipoj9
DUd6urK+i4RTqLzpV5ovJhzlMD1LMriX4NZrO2HHmuWmv9EonXOqJUByTdHS+qeSYlcMZa+isjrtitvtb6YrZC6QYpWWu0DigGENU5YlAUK3V3odZvGMXvx0QfsQBGB6
3+yIaP/o+dGM1wHsK0LNP3h63r3iwSEfrjfuJf8FwQKl28KztJ4g4rB4f0xyQITsvCq1OWrvJGBRAT+RjfdjdTbPlWEY9LyY5vK3BOKIBQettQl/z4WBMy109j8cgoEk
q1b/+EGJ/zXYQ7qhzzstFIVtPZQuPhPo75xU3aJ9Fdn0cz3RZ2BO7k86gcRhQ5L3J7vGQWK9xsMIiQ5bPG2VjjMuivCzH/c9i/dI2kec6fx1TFSs+YMXJ/kHsarbFshM
N/qxjLqWKddxTLb102ftITtqQPU5tL/WF491ZBxdQV4zsirCCYO8Sj6fv90LEABVuLgyiwtKNSpE3ztqSFByn2vuQFyCmKHr2tR+43QTUwr1wFrzLpagZ7mP1ea0zsOs
cCAHdhpqvoUI+XIUSl7I0NDEj869zF5rMBOp/Y5qptPzLJup3x/2Z+xjdyymrXEEMy6K8LMf9z2L90jaR5zp/EMlfMQrboub9l5+bNVKJM7T3uxagNN7U76Qwrkbndx9
ZFP5LMSJ6p2I+LQu3AAsycg20IZVbK+BlhmCvm2P2YtZpdnuTKs8d5c9bTxveqLxGCJrZrSEht2Gae6p0LmaARMjgi3e7ayokV0StapysbDsfDzJsXOvFncz3OD8gFK2
nvnWQrQhkF4LawnoYkDDXNA5DbZKnP5OnKFioljA7n8yPU8GfdaZZ8KjvDOwXJmXNb2rC8dNjwqOq3VQWYrrRZhXYgWtlsgu8ro8e4bg+u402DHj2GVu67H8obR2Cx58
IkfVELHSIBVNfOlc0mt4PinqldxXuNNqhAXfwOGKzMxzVwiM6O31CZZbyfcdee0ejgvPAAWX/VM0ZZ2lG3R1FyNm0GG0G4MVofOr5g8c2wZmJs1gSu+V9A/Lh4GTuQo4
wQtUy8+/khf2Rwj+oR3yz4FAjEi0APsS4jQLeeuAzhNIhDGltvK8HxJd6Efv2gkG04Yh8dXsI2rfVRi9qsGnas93E1iK2Rg5qW9s1MCIEUllxEvg6RgOr7FOdpZJG8V+
abYnoqqiyeLQmCh1+kZ6NKKUtjJX7xIzt/IYlNtHrlPPD/DddbiBy53mM7N48kqR1sEJBmo1olU2c+cgQmwZCI0dhmvxg07GBPCCGXibKujhAkyHsyxelN0IZ4+qPnky
9hKeVpE4C5xB5sxNGHepe0g3ZTPo/GDb6GC2Tm7XjWzPJXwLwOB/1DfkW+KgrLrS7xrPNxn6+WFN5/wf+uJjt9T/D8VQa2xvRembTuH6xlfQOQ22Spz+TpyhYqJYwO5/
Mj1PBn3WmWfCo7wzsFyZlzW9qwvHTY8Kjqt1UFmK60WYV2IFrZbILvK6PHuG4PrucH0ZI6hwnm36Pt2qN0Z1Gzma7fhND+RKuhnLl13PxC3GMmG0Of0cdZlrkIHatF4t
Xtz2fFacxULB5FejHsD+IXJw8Vj2iC04fHzP+xUom+ksTdvAlHY/xAZBovEmSokV4e56noWqe6878x/WkGF7FcYmT/I9t28AEMQKvu8I3zTfE7bp5XtvJCXqIyWYdeuz
VPsIWbHInPLStDGDOZXewJdTwTFg8H5Mci/eFkMG9uczLorwsx/3PYv3SNpHnOn8J/vKt+MfNrkePMnQuhlpj9bnmJeps4W2cRlh+LEDPdki2JpSYMOzGQaiwoifveKM
nui8sT+VA9k5h64bIDfhqwByYGJ3rUWxSKRWkqkTXBowzTrMCwPa0nUafh2QBLA2Y4gz3lYKTPehNjO2f8Xq5AW2v5W7aynK31tBAR+N0vbOO/W+AoWdlqwQ69XKMEQZ
Smor3UY+7QCZJ35/3TK9bFvdKl7SLdBLht2AWsuqdcmVHsvLhSewgLQh2wwmfCUIB2HZEyOOESzLCO/grX+HwFJQWBjSUler8k+2z0YbHWjjU0T+C84l1ca6qzoHPdgI
f1/tlftILZmpRqgDdrWgtXGN0OJfQmBAimhSPnneOKpjyecqcRBMXyA1g8GODUpKF6/0hcTD011U8K3mfFVcs4CHuQCdzWveRNOIN3GTeE3QTPo2H8TCVxsVd2aV7V3h
ZiyjotBm5QCO1JGNcEdgwZ0bvupPSkv/bkE9dD0OoHKdG77qT0pL/25BPXQ9DqByBUsdlkP5SAKfpZMCzoYQyKZc+M9UOUQXUsDgslG7YjfTBgwFJgt8O0Hj4tajYn2n
PdVIynKuIt+e9T+6xgeDli4bpnn1vOGAIkJV7M7qZjCkzCLjlvuV1bqcBZjRtfrCNM6Wj9eoiQM114GMqKjqd1ksQYYOjvJwxNJv6qBge9moKiPS84Bp0VXbQbHOsujn
kYlu/hKOsE9a2OWr5LPC4tahykSTHq9dF7DVL6Fev0LArbjOPNLQA/v2SG3tZ+xxmStNuboyGWfPAmvDd7/IkxLG/DBcwarQuPN9FCKTvl+Hz+fUNiPYPj/ZrdwZlEVn
rpMG6Agq3TEi+0r/eiXpAvDxSBM928Dcra7kBW8DH988itVjflNzeuGy32B/rtFJLQjexIzZOH8jJserOoMGLgqyMVJI8FYD8/MbgPnUMAVhXJZIlWLsJs5gUeOsCNTA
jR2Ga/GDTsYE8IIZeJsq6CLxMeo7qPruUPV/ry/uixdEyxMRIf/C6jZ2eMOui4xeMtJdj1mWFoEmpt0uFRtinH3aU2zVoi6NeEvaFm9aHoNgTsjwdF2KiY6PJDarWTQ0
FY00JQfnxxAY6x4AQmk5PL/Se54ev6rE5uIDo+sF8TsjFx0Ha9z0HmDVuE3ChxL8oDgGAkPCjuR1FW73bdq6Jhy++RIaBweXlub12Lfb8wzBxD67H8qbrh50Cv3Ax0qU
jR2Ga/GDTsYE8IIZeJsq6AF9IOg16QjS78sJ/baWpjghlVfZ58pIoUPUdy/hf++9SekZL5RV46SZ5Maez2sj+IA6PllG7pC6+KpWpWFJWSz0bmyKzQWcw1OS9Wzej+xs
iQXZky7CTdw8RB6iJKWVD/wK8Uv2deupdm8CKghvT/uR3YJz8/8GcGypgXZ/yufZyogm0Sa9h4GMq195YwJtiCNTOF4YAvy4etD4Th5UXQ8YImtmtISG3YZp7qnQuZoB
EyOCLd7trKiRXRK1qnKxsOx8PMmxc68WdzPc4PyAUrZwYrblYePNSfkRA8xjNEwoDT0SnYG0f7m+jK/QCA4BcOZFLcpti9YwTyuZ6w2cN45ZdBXCs8dP/J3oRs7Us3Vf
vVGjz6dXmfvlFJ+BYHwinBnpKvaVzIbm8hN3sTCZ02u0NhAichWugI09XzzTt9dWFKIT91+OAq7tgS+dMx1zkz4w1aKN37cO6d8mQ2RMiisQPbs9cKRIA7SzepFqQ+ju
JpD1T+qvSmcVD9G5HDD+o0g3ZTPo/GDb6GC2Tm7XjWzYpkjC435lFWDFDG73lM8gtty79WQH/9I9Hy9d43rGoM0Ioh5xriQaA0iObFE069J3EkF6bXf/Q1hQ/3NbSvci
R5YB16DIL+BmlIXy1Lr7q003UaY76exZlNfyL0EDBXqSLxkN62Gr9dBEMgvWlzOJzadUtIBF0B2/s/ZWogNYtcROWIPqqK6nnXL4mrsDCJO4PWWyVNecFcXmyL/W2w9p
mIAGIjn/PGdMIcjPlCdpB2YmzWBK75X0D8uHgZO5CjirS7faOHFb9uK9d2eKn0Z3/CPte23Q80Y/zA0OahqGY4vv+0sdQ9IRSSIe0MBUl3vgFdd98i1+l6eWkLsbMpto
n9IYV6vjEB6kqtLBtA1RMF0jTNq/7+mPOhcxqOl9genk6PnO8eVVEtT2bb/ZdJtlR02/LLU1v9kNa+r7WNdDeRQvJrTgogs3llCNn7TNXXAcvvkSGgcHl5bm9di32/MM
wcQ+ux/Km64edAr9wMdKlI0dhmvxg07GBPCCGXibKuhH0wUM4rxyYYXT6HRoddj2m0AsTn5+rQ9evV4pRsyDmVvGrG/4U8NNjkxoFeh2kObINtCGVWyvgZYZgr5tj9mL
s7gJf9Efs3ocibLIVWgGIYfc8hoBpc425yOpJpHoAO7b9sq2WyEAh2N8vJ26EW1G5TXCZbT8Re4O7j+txa4erY4wUO+TxBggGcuMQEDz7mdCy9Gg8f2mgM9EIdlXellZ
IwBq10iZIM/CrqecqfS/nlAJpjFDT3T3ou2Do+lHGiRibuDieN6/6YLGJ2h3d8ySqHzNPKFbXzXZt7ICLJ8TNoUcSOx5fHrbjtJMjGeByNfj7GMOExB+Tv9cCsgLpU38
gxLGfCkQr3hrZfNgnxbL1fXGD15CNUN/BzXrTTTM3fu8KrU5au8kYFEBP5GN92N1Ns+VYRj0vJjm8rcE4ogFBzTg7zNGqwif/ZqhS5xndwVMU3+iVrCzojmmii+fBIyD
48k0w/oc6vM0vQOeEZ8OzZuzlKcqq/ao33z3tuzsegLoai4khDy8AXDAdLQw03nHqwhVwb/e/De40UG5D1/88CTeHeVfKtZF2B3fb175B+qWb0KCDRV8cotB8qt/ffRv
Z3TBrz0Ekvlee0y2bVnh/1MKIBKVyAkrgGIGLASNuTxsOdeMw+I51HrmG1xMWvKo8p2FBN7SzPVTGIYvNT+7ZkBhBMKRiZP89llsEaRytrntY2qxssFfWRVg2rVQEikh
dQSLejmdvzXN2gcbT/iePaG+rLl6+Odif71Ku5jry8RwyKzo0TMuY9Mi3ohGUmbTTSzXMwfm5+M6rukFNrRJjr/JxgeolAL/UizfW6+kE+JeA9DIHxHyNAO5j2BZP41v
LnnyuIFaADfuE8o57xH1a/kp5o+BMdhlQJJH6G7HhYWIYvTiLSLn0EG1tfJWZVF85Oj5zvHlVRLU9m2/2XSbZfFDOUYnBKLekUzkTDzhb+jy6Rhr4YafXa4jNmaz4dnU
i47HjZ6yTMODx/3AIi8tqAjJfE0mSSno6th5b/vETl/3gjwI9sHZehpjz/Ksc40scUj0i2Hae11pqgi79bNp0TiqIwqYhcQfZbgda8NDf/oBMyJeBFKQl9oxva6mUGiG
3/wPa/F9QukFUepRPQjCWR9OB8v1iujQN0KPX2NcXwwFeVK6F3xEaz8KmNfDAIMe527jc+H5qYAK/ZTF0gT9aw61fVAJNntVhMRH2AORks41kfYf0d4dLYBQ6x6XH/cP
KEJz4yN1mZce10SR6Kf84cQhvFjVh/zA+6y2OTtlX4q9bB5knS8NkrPhNEnw+/KVxTXX70VLXYaOAvmQvGz6knkGqPZWeudd/3u6j/kMJ1TcBZ6i6oJIMC1+D83QYNKw
EUBb2w6730SNMdVNDLGON4WUpstATUYRi8tIM6Tx2Qqm/pzIGHbaB7ar/JE+rEsQT0wlefM0crjadLws+P5LLB+KLJVcUwGsRQpvvX+SEwa4F9ugvSpTz330Ft+mCLyJ
ZY3jCc4Za5cQEn4yfqqisiTPt8QGrMSzIsGMxSzG3azsHiPfJegRMQsCQvOjGJB41/um3Evq/98zvQCVsQVGIyKY+f8Rhfl1hmvomgVSUIymMrj791JgmoUhtddpwH9H
Nkil7X0vRYhRvGwLdOQN5j+thMJOuRNnVJiVlP/smO0hEhABh3CXyclOK5e/h1IIeRgVYUzmySosAwckCRh3XuX6qmlx4mlSmmaWz//R6dXqEK0G5GeRq8MXIxsTaLMo
K2XxXHeoibXpdihEW+nfCGcFmkOHgHXAnDYtBwcWe+TQTPo2H8TCVxsVd2aV7V3hhLlFGILgLuNw1yGmw2Tq2QBItradr0oOa0sgsoCZ5bPRpKcS1pY3Z+HfsVVOyFRg
3+G0xOH6C97ml07lcpiiFmQyP3j1zkF/z17s7fO79/C0Wqusis21+3PeNr1m8tO+vw5n5kYj5AY20vM/CPL2UrIt8NRcSNLl8Oc+zxWFYU2JXJx7lMybCFm9HPx7HHJt
bFL6l5zAUkOyfKeNRquqVtrbkL70n/ykx+keJVlwNZgoufTg3Mv8vrsjQrWDU1uv0izTuE35N/nJ6u3OifbZUtXt0mLYoQy/N8XDYYDJt4lMq9709R9PRc4e1SdLT+Ak
wluexQF3+uRK1x+gK0Weaww4vcZEFD1VOfVCZg9a00MQMEg2OMtknADg7Wk+SlG0ZFcSQGNEcBW2AZPUF9uyA7iO7YFLEDkQY8C+RHYzYtwxNMvV6EyrLu8t4/X6N6rj
g5jmwBpaGNdrA0OiaLi1IY/khx3kDJf2uH/aLqZZrFWn7G2L1+gBl8Fn5NwW8MjaW3grrcM/dVqct6MFyjLB8pDIIBdFr9QVBeAN3vnWuZ1ukzbnnV/gL3jyctwZTE2P
7jXM8S81+47Zk6+5Njb114guIrsQd7sNPgmzPZ4Otqmmn0cKprhUz77svt3sOLb40G928hAhXVFrkjFWsgHPMevKNJghf49WPkwmsLvlvU0Jm8zxMW4UKQIE0Yv0qo8g
c7EWfKPAALBKQ/pwuntz0g6mNC2pz6XkP2w9RrBccZabQCxOfn6tD169XilGzIOZW8asb/hTw02OTGgV6HaQ5sg20IZVbK+BlhmCvm2P2YuzuAl/0R+zehyJsshVaAYh
h9zyGgGlzjbnI6kmkegA7tv2yrZbIQCHY3y8nboRbUbNkeXgUbEheOE4Y9lXp8AI/ArxS/Z166l2bwIqCG9P+/x9mMKvedMQj9rdBINon5tzBR9AZ00Ol/vEHvPFTqWy
2bvyni6QJfRdlGFoMI7h8mRXEkBjRHAVtgGT1BfbsgO68hunBlcw4ZUr9m94AtWKi+/7Sx1D0hFJIh7QwFSXe4vv+0sdQ9IRSSIe0MBUl3vgFdd98i1+l6eWkLsbMpto
1I6V8jnYIbl89+tZnk13GYDJMdj/C9ee8xdyMLay8Eyh3Ag2DoV0t7XfZRaxi8pY+J4wzL/hcfXsK+z310otLpWlUrHciYtell3CmWzYInexZ06IsTT81TB0TxpIVPic
QoSpX7Z0LrJOhU+mX04tFovNy9In3jofGt17IIdGvo8xRv6TX0l9noauc3UJsw0hgUCMSLQA+xLiNAt564DOE0iEMaW28rwfEl3oR+/aCQYPTyoJTVJPq8RpdZ0SSmoA
A/uaTA8gL3K5e1UVAzdH0h5kgQczDlhYZoIIsxo8tHsjkJckK6MqAlTAOsehy0QkW8asb/hTw02OTGgV6HaQ5sg20IZVbK+BlhmCvm2P2YuwohNIbxZhRToKrovI6qEk
VbaxSosgazk9RL7CFZzCvNF6ht5rhXlZbCLyuX8nGLFUSJ01uI6Uig82egjM9cKn+/yQLvR0UZNxDMuTor6y1xJWJwSvmoCHLk3VHfV9G+FHje1+2HAexoXoEQ7gQK+u
BfHKrlqMjn2lCcHNCbhNGPsXyNhLpIwaWP78YxfvCPw2WSeHTTn+dGRGsO4dwKSJs+rOB76DbYGn50lpAm8GwFK3BJgpWT/bhvqrFVsWdpvReobea4V5WWwi8rl/Jxix
o742q23jVCFaaci36M5ewc69D6VBaxhyBCpZ9P1MhBsSa7gKuCL5lVHrflni6e0qcnvph7KfFfzmTul9tkE9Hh1nvnIpgiOC6AMbjj/rccbKiCbRJr2HgYyrX3ljAm2I
Q5qFKSByrQma90XlEzQmRzadkHxd+AToQGA5G6FxdN4lALfx/UklBgBv0bODmdcwAcTvF8gwooMKmKArv5m08AHE7xfIMKKDCpigK7+ZtPB310Ecyq+YeHb8SZa3FLc0
VEdLnnIIBWrOydAj13KuzYz12UCPXqZgYgjz/y33OM8Ecxa1No4v7XV4scbYP7pRsNuw7HlOLA9+wkyOg+t7+Ry++RIaBweXlub12Lfb8ww+E36sc9X92iyRdLOmV0KP
Mot5vzlZLFfUdn/rRIwLgnS9qDhVoupG5AW33B4WFEmevIdPkTSmiLJL+/m/8p0qiZzs37mvSCyI+ckyEflsWu5wK0WRUGAHTZNagO81v/QPUTYwe4Tk2b9MtTyZ0M87
HOaP09O5VWgYAxVKywnXWKnALhgyBd1fTwjMvxfX0pjB7qpNqrw3Juv7bVizxrGMMAc+0Pclzjt5fVmuxiYoAg4f/CFPTr7WgguccMNPbHqS5isU+Vq6f+r3fP4Oz6Vz
8yybqd8f9mfsY3cspq1xBEC3OuEtRlEDQsaune+zdB78VKwurpXEFbGzkehesoYRFZHad9pjCXxMfj28uNi5zGwL8v9zeG3Sx107Q3bLQxEXrbrDrX082SM4XOpdbbZx
iJGvWO+90B9G/+k2z3vS8v970MMqfDIrerwDWztThaaHaVMEtyhF7CKsBo02vs0U/ArxS/Z166l2bwIqCG9P+6r7J4lj9GSYzu13+j0hZTLbJArUdR8YYs1wpfBBnOqm
kh/uduzxuW+yesHjim+5x9n2AInLu3P5h7PofnkIkWNpic3X1D8Y6DfauWxXPUkGgO06ic8ZRE0T/IRNcbpRUVHoOAUOhxHhan36sQaGOzSLmwQkOyNIbKzPAJcxrWQu
1Cw7RxJc4RAD+QSJoQtHNZ5A3N7LUk5HO+yWCUAR91EVxXbHaM/eHh5B/25CWXlHMtJdj1mWFoEmpt0uFRtinH3aU2zVoi6NeEvaFm9aHoMco/Z4aZqkHxUB9UyR9tmb
okTgIw7mpEX8n7f6phk5naIOF78Zq9TTEp8sh4mkml9C2fsSpXMR1cdDDkge6uVAqv+i9jFXeiOtuvnPG4O4dIgIP3asJJWTeYkCBaKL4qMvXikKOGu0nWCjJpv4rzDn
4BTjdTLtWNN0Q08c4ji/6x3Rc1kLbccRh9sdeAGQf2gZ/8MVhJSRx42Ku4vV01vHHL75EhoHB5eW5vXYt9vzDD4Tfqxz1f3aLJF0s6ZXQo8UZ3Wtfln1G8rpOEcRooOE
Dhup/zH6Ejydi0L70CGBxfpjc/+BNbQR15UaoDwaJT8nxjvJBVLIPQFqTRy5FDVGGmGHv6dtPB79AeLOGkNDZwPgBUPprdReA60oDfwktCWXoRqwKpFT/vty/DSZA/eR
cX35rYbkWYIip1A+Cwj7WAaCM3Cr9TfcWNF43xl6M6VStwSYKVk/24b6qxVbFnabD08qCU1ST6vEaXWdEkpqAG9ERnuW5YyZDU38/FyznVOO3nkPwdAHnYOY/l5rpg+r
gvX8ZlStviHs6MFUInEaFhCXt7Ote3gTzPOGcx7ET12YcvadVb+2/BwiuHMRDZYrNWKDwlPI2m2uO4HswzIiBZLXjJPB0FEZR/XgvPdc4VTh9d8mMBCybc1RdhtYuM66
dtKGCApICYJGwxmelEZAaLOOMOaXneg03hpnt+X4SMOpGEpTxYo2R2erw7jqlPN6TOmSZbIBzSUd9MvhBCQi4WsSRBWeWND6OgmGcQa/Lk6pgyA+o4GPV4NmlYaCcS59
cNK2I2HVs1XiNv6v3hyWkCTC3YVy81lJ6OzZiYwMa8Hy4eJysbIbOjNe3ntfs4gw65R6iFrXIoqis+xGEBGMh+jB7wWP/TdDfYhyVosSru7DRPqyyrjWKX0FLBqCz8yW
Vr6exgJAGFkO20853jST00CT+/5DYNBkWA22EuCYDRYVkdp32mMJfEx+Pby42LnM6B9zILaAiD0Se66hXXJs8lbysDbc1MW33Z0ITMytC3kzs/NZ2+cz2FVJeJIVy6Ng
EyOCLd7trKiRXRK1qnKxsPSoi7wjo6B5t3ke/kojJh+m/IzCq2vEbpP3CECxj12JBL8a0kfpfKp8t63tw3CKC/3r+1iPsNBcBcPQsmLEiUQD1No5JUAGUlbAoo1RtoTu
WEWsLXPtqX6DrUtJIBT0hxVWQeR7jlqOcm3AJWF3reqfIUvvNH3vdI8vNrnVDo0PI2OhgGIGS87TVsdwhUTzPvjAxnr7PZM2y4DRRFKTQkCONz7VJ2oUsZFkzubQB/8U
+ykrR8RLKstiVDHXnkgXY+WsMn6kSKaFuI91XASjOFFrziP56jEcYIQ+r4tiBBdEn0K9ivdKILXDPltiuZR+KLQr7KJN2JKRMvyprqky5Tlf0JA1ypW4RKCIrdTCYr66
qX35yY/+oWnzEBjcixj2E1jxHwu7tTvwG46Lo5oYHB9E5oz7mr8WaAQoYelx5W2L4D8J2t49waY6rcptutPgHz1QWVoug0xMfApyS4ZZavcghU/B6UHcHM7jj9MB8blz
ynABcufwcDvjK4jpFBqKuB7dlVqSMd6qEgqigNB7C1Bc87IOTcgLSaToZt+lYHjUVQsuGOdS/sjwL8ZOLeCGEd/ACfj9ozEqcYLb2L5HC1+OMFDvk8QYIBnLjEBA8+5n
yuHp0TyyjnvblIeLc1sLW/D578Ej6qRi8/n1coSdswn/ALDxn0rDA2liWlB5d7+//CqeU2FA5UKtJgQccXsxjcpwAXLn8HA74yuI6RQairjvTGr0a+7EolDPLjkFW/es
8+GjWdIniZJA4xKYikKPphev9IXEw9NdVPCt5nxVXLMbnTFKTrxL4l/qQ7zbGxZJy4UVwXOvgYT4TJJsqckut55A3N7LUk5HO+yWCUAR91EVxXbHaM/eHh5B/25CWXlH
MtJdj1mWFoEmpt0uFRtinH3aU2zVoi6NeEvaFm9aHoP4Q3gZX/vZcXcea0htz1wxCAiP+UK5pBgU0GD1afyYrWJXDGWvorI67Yrb7W+mK2QAcmBid61FsUikVpKpE1wa
MM06zAsD2tJ1Gn4dkASwNmfOZaW12eyq/2tF6Y/OJnHNCKIeca4kGgNIjmxRNOvSdxJBem13/0NYUP9zW0r3IkeWAdegyC/gZpSF8tS6+6tHzuQU33wl9HYZRHomD62O
mRCghOMXlK0EqPEiFvlJh/a/EJyyR6J2iuSBYMPqiN+FxSd4a5UclWcsZW5itsQma5uw0zKSKPyKbbtnANAx0LTPTrLGggoiiY0dpwEMNLMuyXSvTip8KH1nBmbwpTmx
TjB0E4D/XI2NHc+EJmIVI4j+41bml+OhWPwdisz+wZotCN7EjNk4fyMmx6s6gwYuCrIxUkjwVgPz8xuA+dQwBUeJgouMqnX+2I9/CuZ4cKBtYxEnDBItmEgkxVMpGnCz
IkfVELHSIBVNfOlc0mt4PhizFqZXqyHg4KEi5DZ4OO4KWAbPbGDUabX1pCYH5Mb8QqyhZjOev+mdwujnuci+op8FmiTCF90lCl9I+aAv4YHb6Imtr0S+AdDTkldK+5Ei
uWKdhCv3F/3QfksuiIDJeuk7LMts7H02Csu9g6ScKZ2Z+kR17CuHFkzYOA/tjEYIqo8zVTDYJ7PG2HH1p4Q/2/etSo46JNIh2FMgyDkdWK7Q87KD7qYVpD8a8dgROe3a
jgvPAAWX/VM0ZZ2lG3R1F/qvQibmiZcgwZP+ORhydyq8GzydFyEBIpxohBFzZAJbwgwYG6feZTxrLgARj0ks7JkpmFdiklxoNTKgJiSuo0Qnu8ZBYr3GwwiJDls8bZWO
HHsev11IUqi5JfmWkQiEYMgJrI8vrHkThQitU/zEHauW+ccF8F+I/ICJ8UX8WV2BpUqcmoALovbsDvDHEAw5xtdjZlwkEumFTQKVPRiPUgDRd7jwieON+SbFytAlsXue
zLTfg+0ftuVBLja0AyIbJ49NiLyQQzbOw9EVKinOmuIbnTFKTrxL4l/qQ7zbGxZJCtvK9uuzNVo4Z/Eo9iM/So2EEhe9DHI1QLmvfYTFZo+Ku+t8sbYADGua3ezHvns9
AraCG6rOiVuo0XAAE3BMHpsCw5rBhLpEXizu2dq1L+biu/bGdLM72vejoedP9x93i+/7Sx1D0hFJIh7QwFSXe+AV133yLX6Xp5aQuxsym2hD26jdEA56MPvI+QWsjXBl
BHNrwU1YIMyjceagZwK22BeSbJJagDBnAtTbuWy7fYWbQCxOfn6tD169XilGzIOZW8asb/hTw02OTGgV6HaQ5sg20IZVbK+BlhmCvm2P2YuwohNIbxZhRToKrovI6qEk
VbaxSosgazk9RL7CFZzCvBhrL8i5SYNsYvVZH5Strzvd4eF/LVKWzCWBhAZ9Fq4YqTZSR41bGPSAKZMXcghUIMpwAXLn8HA74yuI6RQairge3ZVakjHeqhIKooDQewtQ
XPOyDk3IC0mk6GbfpWB41IzwPk1ZzNpUfY4v+1ezqc/hx2marrC1jGznf89XTIGXFkuIuzbFohy7owv/9ddN2Fzzsg5NyAtJpOhm36VgeNSM8D5NWczaVH2OL/tXs6nP
4cdpmq6wtYxs53/PV0yBl7Pqzge+g22Bp+dJaQJvBsD1V7kYqIesltROkhqgfSPZ8N1aPxmevwymdDSlfwHvUOWsMn6kSKaFuI91XASjOFH/wKSrPxJRV9gDJH236QM9
hB4TeAMDFwF4pDTHRZWvnGm3KphmfE7yWT/9FwcvcjuK80IToUXh6Vy+ChxB2NJZTd2Fl0IrZC6n5HJ2RksCZfnCJIOwryYeh5T93mEMESIySUoJKujQw6bLOIdp3MKi
mLSq2XctITM6bb2bNi4WZStwd3R28K5kzTUlhibC9NFE5oz7mr8WaAQoYelx5W2LmWzqLU7ZNpBsHGjFlceyu/8AsPGfSsMDaWJaUHl3v7/mPcKH2KFNHq+h1K7cIZ0a
vblKj/Nq2O0/2ZerRTEmWJwufKdcN4a9SKCKT3pQoH8s0h1GzjAR5sE/sJ4Eg2t5DyFdKloitTgvNU7qgsI9OgEVOkucnk0jxa57iHwJ+gdbYvurr/0Nl1DEnXE4baCr
8yybqd8f9mfsY3cspq1xBBx7Hr9dSFKouSX5lpEIhGDICayPL6x5E4UIrVP8xB2rMTweFJRzWBJFOK1uCVsovywTQNkXIbleLNRvcLmk2b/E+6JTOboFZ6ue6TB52Wuu
BqNtSSmMDBJiwKY0/NaMCrGG2vwPSobZLIl55lrmAtTkPOfXWTQ+q1c1n7X9cvHHfrzYUWlSpFYu7jMHdgF/BFm8UG9py/HhKGFeaDxM36CyReIFVhlfQSI9A+vra32q
xGqK05o4qouWhxycoRjGmGQBMTVrTfsecvg04x/CQdZycPFY9ogtOHx8z/sVKJvp3z4zXTHV+ebMNalaXAGav2QgnU1EWf/ntKjHckrqMU0mZZkTO4S9xQJ87YnwmYB+
WXQVwrPHT/yd6EbO1LN1X5gcI7XgxjbUQDjjb4z1hVVE+s3cOfadoaooFicH+0tNcdu+82m1z1cgCeoKk6iucU06fK3pfHj5b95JM/gpXMO3uxC1G/9rDclBDv6hd8xw
D8Qp3FP0NXUM7stcjcVQLcCtfuOZiSyfGCmxh0ML2kLJatMs5YEpHGpo7spmx2O80t6izK91Exnx4jMXkrHLqprYDPmjxKtQpbzApNKmhVw43XCnfG/JJZSXxQkmXsLv
dBGFIZ/B8/PSaGXoVzRMOm7WMBnGQJ/PLbqb1cDRA2nW7L1s/kibgvQjbjnrW00tLhiuw7JB1l5q6olhxnKNugcUCaTsG/rFXTB+eBSUyvhL8PLAncC21WNfxBbOdyb2
8ysDNvmPpUDmZNqAt6794N/fa8/f0H+lKui7u9KiBqnsW4ncTdUXdMfvDqp6u+okidwI05hLqiDKYxBLPUdZIgRK5jENRLQru9h+NUtAAj1LRqvNRVP9+LrLjU9YPSU4
J9zXX+2DdQLngUsutO2muGYXls3ucJNqkdlN4lesRy51W0PVbQbZlDtrI/NUn+JQkj0WNWoT3H0h+YGM5T9hrHWSudaSZ4RiQVXE4jIHnrvOaEdiNitYss7kQelk9ERe
0JXOuAfjBVPacW5dF0Z0MDxeB7bhnvsWJJ57+wA7sxQJbG0KKE6xQ/qE5+QMsaFMBknZx++h2Lpkf8g1Y1wmNJOwbEpCP2BEgneaK5vA67ba3i0q38Uy5r1I3TvGApI/
Vb6lPFBM+l5myLBA93sZO1ml2e5Mqzx3lz1tPG96ovEXPhYNh7LZHrruCWqyFvDgzVBZPCYUjFwMnZXtmmlcs1Ak+2UauCu9xfK7PWdNkdSZkgOxWfd5V3FNJN0Yv3jA
HlwavH9uV+uFB9PIp2u3HqPMIbOmAVtqf521RGW3OoVNFDo7Mztuxgq+UvLj8dEIM4x3oj4XPPBehzDSjf2sAI0dhmvxg07GBPCCGXibKuhWWT63iQKrWEnFBTZ76V5Z
2t4tKt/FMua9SN07xgKSP6vldsmLaKN/DXy6qUqg7D3PK0R6AscDAG5YPtPI/DzeYhPe3nhq/WxPqcMwrrOSV2g0WNHs/JFCbCbTb7DQu2SBea7hXtw2meTe6cRdAKBh
vOwagk7Hf/tIcYs4ulgVvaKly3HS6XmiGCrQGDUfwCXh7nqehap7rzvzH9aQYXsVwLDIndM8JiZqHxjQ8vDYRiDuvmhJlY+jbCHJffOinjv2nmDMlkdfZ7f9RxGORBza
dlr3X23/4z1ZHzpD9EC1vjrtfBkjjqBlKeO3kxJ5+E8zPPzHWtnf3OQhSyRuWEvPm03TjqFAc8KBuGUSe3pWlStC6xtdlWwboOH+eJU2av1B9sBH2BTqStZiK3KkylDC
xIcglkxfoAyX3ug90OLDE8KNn6GjC4C3MEA5YiNOc9HN0JY6zzHi9YMgxzITlbgjMzz8x1rZ39zkIUskblhLz9O37In3uNtzac2k/H60wDGRvvbjlrdVWcXr4r5Ex6sY
r7mIDdDxOOP3OF3VQ50f7bMJXxI+011rqWjcv0qEb0YFKzm8p2QJKuBnpAIdfKem6/GEA6eWSGAjlxwV916vQCFP5sUW5ulFIsu5BKF59EBhBp55GLFtBZcSH0ax27HK
qjJqYyDySnealSXY4HKV/raoZiZXg7Qu6Vg4CkhAQSipsymwChi7rENQpnL3eVYCtqhmJleDtC7pWDgKSEBBKGm2J6Kqosni0JgodfpGejTn1a3tVwySU+RGzkG8dtsR
8L4skYJXdPy5d1JpfIMmtuznsuzbnFMZMFnRXAt33SbMtmLf89xBmUwjJ7TJEzPfPFvdYn+A0LbZq3ahQ7jCAptN046hQHPCgbhlEnt6VpXyEpNU2/pvuntmpWYU0TSO
qjtxLtRi/Ioi8/vcnhOhig/2svE3JJHxjN0Y9BrXDD9Yya3KjOTeakFinbj9OkDhudlTxSBLJND4tBxzymrazyOO1mt1d00lna6BufqK2DhP5j+90Z30Xc4nxq+xd40E
NdfdW9I2w/VYvdP9Ix11qqrPkJnwOYFaowDysCfSAUsrltICWRb4i2yEaGMMT4a/qqPtG4Pwp1kVNmuR7XNVH17HFpnk9tD00TRezE/9rFatCAk5f1AR3S4W53dXKrZj
K6NcQ9Dk+tG9X3eUofAEiUu/J8KlcNjUBQ+hiUhwuAOpy36rCF5tkwVG6hiFcYyNUF6AGWIK2T9zx5IbYcbM5+3C9LteEdzxuDFakgVLeq6ZC2ZW6RdUdG5n6EhKsMmd
bcOQHoztWV4rdB0wvaLP3Xdpmv59KuTJ0MQUlIQVA/L4jmC3cC/kM54/XuyJJKlJUdJj1X6H4YT98mpdABVdcV3qvix6lkgCSwtMfTlvQbBNB0Wihh7WpYgySPpnPzPP
UF6AGWIK2T9zx5IbYcbM58omU9+MzuOXvGdaQjY+WFCZC2ZW6RdUdG5n6EhKsMmdbQwGudRn1hjjpPbAFxfPvqm7qp1+U+4g7nYhby5AbGD4jmC3cC/kM54/XuyJJKlJ
aQb2b8LHhiycw/wW5ok4aq6kDyDGR0KniNSQrnUOBWL9WgRXXXTHOvnT193KtXIxqACT3qe/KtM9ki2/WcbtQWKsRJssSxl3gfDFDMEse6hNhR97Sl7e1hfn4KcwJ1k1
hvagvtNP6UXnqstv6hpiWaKXEq5qj1smwcAU8AqIa9lexxaZ5PbQ9NE0XsxP/axWev5x6tnqoF/vHgSO8tM3DnkGqPZWeudd/3u6j/kMJ1TbGpFoyY04lJW4eBPJ9IAg
abYnoqqiyeLQmCh1+kZ6NOfVre1XDJJT5EbOQbx22xHwviyRgld0/Ll3Uml8gya27Oey7NucUxkwWdFcC3fdJmo3C4ePAtzGEEqa2gAgklpDAcjHZlewUHya4sKTAMva
ujAVlYcd/usgmqpTzhfntxk9Fw5IFnGgrEEGdpv10nhqNwuHjwLcxhBKmtoAIJJa2Gz+6+mtdnK9+JGZyHmx4WGDG4yYICz0LXz3owc46xqhUMck6S0Ms5pjnRt6961A
ajcLh48C3MYQSpraACCSWrSIN1h4JhWR4HcN40+oTASUTzOQPzSOFiCayk6RbtjMvO+uWuJcezn1lG0BpnP2TouAbcVumgfMm0lRxQdxnSSfmoTo7Fmjfn7InDWkpY5C
LrDME2sRAJu5CtYzIA1widb8WZr79VvPbUHS2C+VDgJmn7ZMHcrl5bT7pgLWUvpiioo+taTh3JYX6kPP7c+ZBDExCx77eAE4ckr6y2rNzlR3EkF6bXf/Q1hQ/3NbSvci
QUtnLG4AoaUkfM0gK4RNKIGJ+Xn+jwH44t60OANz/kqTaLTQXYQGbvof4ZG/hkRwabYnoqqiyeLQmCh1+kZ6NOfVre1XDJJT5EbOQbx22xHwviyRgld0/Ll3Uml8gya2
7Oey7NucUxkwWdFcC3fdJvAsoxYLLUywyRkFlK/VIlZigoJ8ZtqWUz//Ze6f3GbFi4BtxW6aB8ybSVHFB3GdJJ+ahOjsWaN+fsicNaSljkIusMwTaxEAm7kK1jMgDXCJ
8rm5S3vJqbik67KNQXshup1ZeKvDyRM6NCbALlbWhMGSCxSCiBTQVn5MQLtijmkXgUCMSLQA+xLiNAt564DOE0iEMaW28rwfEl3oR+/aCQYYuSSElke2e74cnSBEp0jc
pj6CqgxxdLa6lDKL0ew241BegBliCtk/c8eSG2HGzOcUohP3X44Cru2BL50zHXOTNZazkW6a9J7+tiqs2ud09sc/wSwgSLAKk6tfjuYlzxWH2plCUoiuXYZpnhFsx1he
yw9H7oehKAEwFGXyK78O350bvupPSkv/bkE9dD0OoHLiX4K4Yksf9F88cX6OtDMujNHer1hFZRM2EmsCPgPJpIDJMdj/C9ee8xdyMLay8EwiR9UQsdIgFU186VzSa3g+
KeqV3Fe402qEBd/A4YrMzCMbS3G9M/fkhJsKBbYBIbHi95sJRobjJTqzFVBiAx52oLquxV+JS0qxKTWMK1ttpQ29cxPJRSqQe5uUICdP5a3q6c4aCTvbp7oEH5O2YNnn
abcqmGZ8TvJZP/0XBy9yO0XfHU9yAvNN1UWTfJPnsU93EkF6bXf/Q1hQ/3NbSvciMwdX53cGL4v80dh8IylIdl498dxcv7I1HnCbStW/MpLp5c1T8lTNTreB6KtRGvZM
Fk8b2/kU6DOHHqYHhq24KdisN04lhwrL626ka1eItIB20oYICkgJgkbDGZ6URkBoBp4qSGAJui63JwX8diYSW1TadfU9lMYnVp3WXCir/IZ3EkF6bXf/Q1hQ/3NbSvci
FoG8Zr5opE4YeSYEbBRHx8Zrds8d0uoejsyYjzg3yzhgw0vi5z5CWUnc2X8hDPT6lxZA28quLa6e0bq0s6HuwHI1duj+L+/LMol/r3MUiabt118pVM2FNN0Ie0Q5KBEO
q4YGURqI2rfDGqmBldxufVsjRrZ4Wtb8qmdhjzBHMpAx+MuKcvD9yxOVDZEUJvOs6EJ9DYRMRl9bBjykBEZK7lX08xnhOrIzOmhBFoXE64MBXgaIPbRvR4O9HdPeJeP/
m9LeSvpJxfm4Q12rB3cPtIy1O2oYsXwpnq2MFvYg2ehDbLsiCZ/3pFrdiZtYn/fr6skv4CoQi13uPMsJjuWcX7704PDOydjr2m4bz3eX+jgVNjp6yoz2XXss8mVsNuWe
WxQ69LX5T8K1M8WRkw272+cs/DcHhEZhbx7eAUHN2v5vKbOeAsxbqKCOf4IzOd5zxudK35mYNkFIyqbTx1eJIBXEFWDU2FFNJ24SFDFHPrOplHO/oimgxfmeiuRceW1q
Gc3uNeCMbdJwHNWEszPmMK4l84+5A1s4PbMPENnv/lTg8T7p8s4kLrsYI50TXqkxyRdjfqv3N57F6tBDEwXeFQXIYpmNTz2luAXWIcSHT1NruJp0Daj0EnWfgQHTetrM
nwWaJMIX3SUKX0j5oC/hgZzSkPzwwl+CKkFiwfBZMHDbNN+/JKn5mpCDuRztLtcf1U6Zaij4gVF0fTqKWIEzzVz2df8Ge7RETjXbSs6GujBkm4p3iCz1r0ZcXhAYGwo2
9HM90WdgTu5POoHEYUOS93to3MFSbnzkK4O2D6F98DqdG77qT0pL/25BPXQ9DqByAcTvF8gwooMKmKArv5m08ILHA7QoM3lJa2GJgTg9F1ZEclTwTzUD0V0n8e5wdhyz
gscDtCgzeUlrYYmBOD0XVr+yyBjnLJW4hLOzy86bgo7a01OMvUgj85a8yB0W3/HoUB923LDMT0rg/hltxGeE1EH6RA6h8MQUprdkcVRN7vwg7r5oSZWPo2whyX3zop47
6I1klSFGy4x7yI8ox7w7Y3cSQXptd/9DWFD/c1tK9yK4GvGK4wnK/1e2MfwCTqx3l2J42Be4xKhgYnZGv5tIDyC5oj7rCf7nzgAqVLTTfVyM0d6vWEVlEzYSawI+A8mk
XPOyDk3IC0mk6GbfpWB41KzOCncb0FoATAp/LYTAlIdguOWBWG4i/0huKnzvh77ZnRu+6k9KS/9uQT10PQ6gcvx9mMKvedMQj9rdBINon5tzBR9AZ00Ol/vEHvPFTqWy
xtj0hFdAfbpgN/m/yYLUXj9cRETf2QB00lfVcgqZA2N6tox6npPn6JB41lj0ozK7/2lkXqi49QKS1TzA2boiDhE7wbcMYZPcBMlCeRp2j9T1czva2+1EePY9fGQHSuY2
hR0eQtSVhi60CM/eSxNiJRR6fJQK7eiMr6xfU3uvj7TMtdynicCyGzqFl0ujZqE9R87kFN98JfR2GUR6Jg+tjmSFNGOwCF8fw1Hi7Sf8xmuqiq3WEdnEpA52Lhw5PbJT
X5LzblxKFntS4QlS+3KvYDLyL5SjU32GDAOtHRVSCXDQFA8XafE26kN9N6ssitP+M5X5+CIBrOqJdsR2+dDCGvLusni0wiOLhqUgSEI/wp4TENmOHrHrJsReWqL1TEml
pMwi45b7ldW6nAWY0bX6wqqKrdYR2cSkDnYuHDk9slPf0mROK34wROX6dKy+ahB/yneuEXwIGVlHvx0IUZw1lNaGirY4JpF05HLnSVDo/HedG77qT0pL/25BPXQ9DqBy
3xO26eV7byQl6iMlmHXrs1T7CFmxyJzy0rQxgzmV3sCXU8ExYPB+THIv3hZDBvbnj871AA8yVnKBfd/LfycH3ob6zmZ9zQ6SnSFZxkvWmQnG+6H1YgD2YqnOqQvY3hub
f1gY+uqh3hY0w5c+xQKxLfetSo46JNIh2FMgyDkdWK5cyGRGBIXGpmRYhKtYA4JJR43tfthwHsaF6BEO4ECvrpSZv2VWo4FeFk7AvITjDlqO0LwqeDPQGMrsVYhh4lR8
FERtjrwiz9ROp2BU7Hj+VgVLHZZD+UgCn6WTAs6GEMjlTQB9mldjqx8tqq0rmNH7MPsyIABBvKXhUfFzQ4Yw323x6kOtwsmNMT1/mE8imOX3LX6kFkzfgM/G6zN3ugy2
1LZBiO1W9YgstlmRf96JXsrvtEHogS2pU5DYQ0Eey3FQHiRHLVlhBiR1eq4jFf2I4KU8pRiQYkY29hI3F7dMlCRAUtuOsajKEq5OOYsSKYWVpVJSiDNGJk3Fwat5o3sY
3A/PxgQYWgYJCytdn1VqUeHrwKPw3HcAMvfJgmyYZF74n2H4qi8YEwJhBr8yPk73kmPctTsKh7jQAG1hvj+fw6IpeR9yKSRAK47hVCNgOnROuLbAoyya9CITBKgC3W/y
qLoAk6cnzTLBHSMMTGWx42qfzTFwa4Vv9QwZoeQw0IRzjpGijnySJKGwWpX/GN9GILI0AFpni4MFehUXs/f/Ptn/aKugH1bJJSvfUZIdCjQS6kBrt6uQCHYVzb48YQX+
yweD2azgD80sNl2AvSgxdiUBQUr3bbl+2OzrMNjsbu52Gdncci4JxxP1lPGZ4PlNGv/Prijtm4RWA2wT3GqYYb72+km3WL22ofK2Ui+hwoSyZEimeuCgjky/PqWI7BZJ
+kC3P1BdI7+HcWHJxLIBQzKVI40OtFdp15GOTDduO5HZUBDE4PTEHpCPIxDq/quxllxOG9oyDz/IoF4TC79JEdlQEMTg9MQekI8jEOr+q7GiFfqj9m4r4/+zOFkA7zKa
lxGxaK8zI0pqjQEtofJZhJ02EhXZf3Wlf95jukxpY49Q/KPvhYhqlMFu6hD5lAeGm9gTYeeU0JPm/IMCBezRaTidc7iPpV3COd1HaZU5J97M+LC0ueSFVUeWlUuOCBnh
7mI4I8p/NDLayTUwAX+ArJBQyzSN1B0R/Hgs4NKOyuGgzhyzYF6EQwBip9rulDrFdX+YDlpvYrq3kEsU6NALldkUkRhUpu1xxYYmXZZgJO3SEKPHDZOU7Goma6YiclEw
+J9h+KovGBMCYQa/Mj5O9zs6XGoZw/du6EWnUhX+2DQJ7J17qpAxjDIJxLeYg6u7+qXIvtGzEUMyAaJBlU4uNyx/RPObuapl3VuKDDcTbKoq/y+RaHfotAzhQrZrb6OC
7U+Tdd0N5dSNAz7q9rk+KE2doekEMiIE44X+ge7TOMnD1GnlurMQHk7AVpF+QH19tKTwGhGAMnThi/rRMbVyvdgm4GnRzForVwo1SD/E3rcE6gDCRp+p9kGz5BR4SDGW
sbCxjhTGUxZPG4usDxQ8CNij7cRUaJkY0cV6EHePJT5DCnVb8tXa8vg6Fdh+psABjRAduXOS+JEmCA0Fn1/r48kni9dTZ/9Rficjr+mqWpuBplj7BNYu/ZVrmsO1eY+g
OAxSfXCWYeImrqZZam07jq2wJSltagSoNlNSamNcjm+jL7Xj8oWuLiij6ebfC1u8ifr1Q65EbY4ml3iESOtS9uHpir72V6v9P7IwtXZ+RJNkdX8eWvU7bgZTwe4NG8Pi
beUShdyiax77RzqcZ75g+wg3LPgoRV/dXxuq4t6hNVcY0Lpd69KZh+rnoJwMyDq0WAX0aSq8jdPnfYofg3WoHVrmVc2ehNYetuOfq/QTMrYU5Ihncfw0gatvceOWHAvA
oVUg6+gcBFVkYyJJXiA6R09w0qZiybDf7bbxqkOxgkEdDzvCjNT77i2NpjkAPOm8rxckGLhLTTp91WYCExKPqGSNvujCRsLrRe9Ukc5bPJTl/nhwjT/CZxHFlV6LRSr2
oGMy9b29R90b2cnUqGpl4kqTY94tfXflHzVDXFQZvDvIa+EhhBf2LMNyAUeDOceZr3RCnX+OdOMgbl47rwddSm3EEwdwByVc+Pb5TsR2awXR1g0v/Z/N/4jcSjvUuw0B
8EAXPadTFjc8jC5834fDIv1J5brvpnjOkGpJ0yHo9/2NbQTUdC+Nb8qwYW9drzAobQtC5dbVmEupEXyES0I7QuhSScxuug1YoVAK++T9eO2+/LlEru0AOdVcmjdufJsd
BL266BbwLJv+M4tXkKaf5lr/iDTrdPE7hcrrbuVtONW64GLFTYWXe36KvZ9TQhefpU9jG2s+QQG6k0tM+Gi0pzyrsVybILkFDNMo1UtBKQ+luo3EGcGS1ohZbFYBSTdR
S2XgYDcbwxsURaPm3UQcp69Lgkk3gzprte599LPveP3lTQB9mldjqx8tqq0rmNH7A6/pPhcelTvMzDANMQgQ/2hdcYL38ooJlztKP+I13HCeYWjzdzwhrNDFY1tx3p28
/4BpBgoqA1x6xHxRFn5paiHc1BC6+jhjfAgObw4xWFEW8fNZuIJkLL2opyXzM3W/j5Lt5QUXfdmAVMfWrCc1dN2frUoTqVGuLRCppXr8f7wYjXC4aYWsPE6qRbEm3Gfj
ULCEZ26vvOq+fadVbcJTTCBp8yEWG4dufaL5F6K7Waxq38xPR7XUQkhT4+k0sAnSADzOLRIyu4mLDebjC4CN/FOhCDztSP9zndoGFCBnj5bVHpU8Nsm1MCxTuuLD126+
axDH9gNYIrIvKQGrape+OVOhCDztSP9zndoGFCBnj5Z8ffPCXAY21wyL6/CGuG9uLn2d2Ok9xoyrq4KhlSBP0qLNv/rOC2VRacSIU3LCmLqqeWq1owsgB8D+xRMSWKwb
dtmwfzhChchSh6UlpVdBDmBoZFPV+JOaKUa1f30E68L9UcEXHqW0le1Pgro/A/5owedYTg+t5Z83M+ce19jArtcUKTjbZ1rDb4o8eXLxXcBAJaB6qvFG/vfAM8UpdbJf
3rR8GBKbDIJp+vN+9qM9lc4eaY1bBSOgOk8mVgwbwjH9i3Mq8fhXaP5QQPWD2xkmHFnRz2MQdfLjJI9RJoIdhfXHIv8v4vOReQBrd7wCYQPQKurmGyeU4mxUkwAjeai2
FqL6ozc38Fa18fy2vxZM9+C81MU7LSk+eo+gRNRGFCFQ4UnBkDIrATBm7se0jqV8HE6t1dTGrSYngr6zsHvZiyQJFjHXE8Ye2lTxNm7YeNprjkBAT4K9Fu0Qt/XM+emi
gePjS6mAxWqLD/d47Ciu2cBHGkdCpBEVFc+Y9V217TzhJ/GtpzphEEFLy7/0nBZ98R+mP3ZyN0yhx1hWnZQcSh82vi8OBFHtPcRiBOOrWsAgafMhFhuHbn2i+Reiu1ms
kta/zod0Fd+c3HdXW0dWYlDhScGQMisBMGbux7SOpXzQ5lfpdZziNvOhVjrj3Ma3t2X2bI/12l6Xb2UCIWdAZ+ClPKUYkGJGNvYSNxe3TJS6iDgUcJBNu2vd8W1Wppwh
LqepOsghBfdEizs1RXdqFxCJLOS+HkbD+vejgUAUYcF+FLqUoYWgfB7tzHlVe3fxwLRaLWJA28d8b9WibEE5FRCJLOS+HkbD+vejgUAUYcHiyN43iNeFvHBlmcUGHUm+
oHW4Nmp7AM1aZLDV9z+Oj74kbrPNdmJ+3mjeUC1JXzEyIy9TlPy2ztgdq+JE3IdXZ0yIVGcWE9j7W0WF9Mjpj8AFbbMh+7gGgcPcRriXyTMgafMhFhuHbn2i+Reiu1ms
YU/PBH5kmCDunHKyO4XivGGcnj/EMxZnab03hTROc5prvmfC0bStZKXmrVGhpYpYn4SWfCcpHaRTW4iByHvGBpTxTY9+VSAtep+PYBr1toIWovqjNzfwVrXx/La/Fkz3
KyOTFVIzuSxJBKq4GKR8lb4kbrPNdmJ+3mjeUC1JXzGQl7R1G73J1Kx0A556GbKOXCX+Y1hYBk43810Ah6XrOdkUkRhUpu1xxYYmXZZgJO3DkAzmmhyBCyjvci+KYRdX
U5sfrIsuBQu+vYP36m19UN2frUoTqVGuLRCppXr8f7xzOiHGZV6fLwKbnZqpEGRoFmh1SCrGplxZGeIjos1KJ+trHVCQRpp8CAK4u893V2PmPfjyEy7amfEfwLzfap3Q
6Q8BBGb8j46oeCkjVW0gqCBp8yEWG4dufaL5F6K7Waw10f2AnGuu9NNtS+zDlCAF6ZWQQmvWXfgbUzqMqR2pwTNv3tUF7Lk18y4HTUBrwiOnPIGFr0uuORr0RJs95N3K
2BgpzMpqo3IiCSMNPNRaLxRiwHZJEJ1ypqqKgExMB/Yjqv2FPP3F4EHGoI81CzUVNb7jMa1DC8rVfuLdEGMRAkYJvE+Y+H7SN2Ct2sZ0flMGluUryr2J4+dg1RDib7NC
8MPA4ubUgGWZFGbZHApNOtILvtLImYKbqdQNjKCXwWWnPIGFr0uuORr0RJs95N3Kln1o+ySC0gNmnM7SLHWdEetrHVCQRpp8CAK4u893V2O13iyXI5iNjGcw/vTnaew6
FanwuiCjeVVA/aclYudD4RxZ0c9jEHXy4ySPUSaCHYVE29D3JHGskxIUD2MWuBHw1dD1b9VINxG/TS/mRDLCjZn/k5JGhhcK1qY7zmqqg+U3hEfvCi6ZyB46WjTaVYj+
ZV9mk+eOaZc7ibLsH5KKjhudMUpOvEviX+pDvNsbFkmUt0nv+3wc5i5ywIcdPB9rHQ87wozU++4tjaY5ADzpvPEyQAqror2nUj3rXIObAI45a39oVwlTdcxCW7tiDXVM
LRz8ND7Ll3bRTID1h8apj8qIJtEmvYeBjKtfeWMCbYgmmYL/64CSWoELjaVWhKI7U71lmNBrB4z0ucHALQfwNL9CpZAzvVe0vjim57KfkwROMvncwnsAc5jOzFmp+42B
02LnP244d6bJrYgd90CZ1GPUhFXaI8kSKykRqOiTYuMZzFHm90LY4lAHVEjoXGg0te8Xt3IvuLzTgy0/jbTQG6J3ie7uWSP/GVt/BENsUaMI2W5xTqJY+oHgKesws/ER
GY4+rg5G4K95rFxsT/hBUYYluLLEEGAVohtnPTpae8c3YhJGYZiy9uc0HbPA9G6e0fb3+6yAsDEI6uYbAqtyHax+Dwn61x96pT1+Ph6AY7BszlhJys5+k6/hcntH6M29
K6Kh2pKDJiA4Rsm5wbL3xypW76ATzUVGV+BXDgyZHvCCMhj4bx5No1I/FG48RbgenJ/ke6EXREq9YL0GI/SkXORooizcGhpQhOhi8L4Z2nhKXLjPRLG2fDRU+2fg0hra
Dw83KT8OBSlDDlzximYIzja/tYFMH3UPQAQsqZqxTIzsAF300tmjyI+L2k444QJ2i1LfSHL7meCZLO9MHcLDPMrLTBckGp8lwUhpGaNl3wAfuqyez7d2uhs6v7M6pAhb
oF0WLpz/09rXfCGzxsES7tcUKTjbZ1rDb4o8eXLxXcDK1gN+edQTPY8i0W/+b+lC0ZV2xJ0BbMzywXVyUIrkTaXzf/oxGPe4ao2W2PYTFf/Xe6rYn7oZDyG9/PZa7PSc
WabCSr1MT8trU/RcrHT/1sK+JfPX8kyjku0sIqXdcvyh8VTo37hyWY/SlyM5cg7A6C8LdHYYunW5LOPuJXoDdGdMiFRnFhPY+1tFhfTI6Y+ClYaabgh92mQOaX9SPnis
iKGO5j7T5NM4UsabZgPjZNQGJQXfl7N1SoJ42fFrCv2Awy3rOCbClCBUYlP8RG1QJyIJ/TwHcVIxkrGwbrBPkx+6rJ7Pt3a6Gzq/szqkCFs2TwW+j1N4fOyIQzoPZ1lP
1xQpONtnWsNvijx5cvFdwAbqsEYQXLw6yNZHOVLIuknxgo6S2FjIiZAxtGi+DwOZ4YUId71VqluCPXHi4DPMmGrwLl64OawgpciVwHHnB3iHeD7qaG3dW+dRWzPynzpA
nNyrjjaPlzOJlldz5Pc6NbuZgVie1oI/A0ys1mmCdtoBYpUlBInpWpnJxKzzpAK+D4uqU8s8r+u2h+dwxlFyeAP2vGydxVmE+N/1DohvD6OxLJToS4d3h5hJ/sWUhKhT
ar1CBOhMVPvMpmQoRzSxKoER52Sh+57jqdg+0kNYWfYm24XspQBKtGNsxl7BgwojRNvQ9yRxrJMSFA9jFrgR8NSLgDWUDUOdEkcK42aDtaawSwdvc19Ms5z8BMRho8Rq
Iz5UyXPmhOz0s67qs7RcZnrsKz9QWesrwTEUYV+HGNScn+R7oRdESr1gvQYj9KRc8xAgFg5xXGFwwtqipQwWGiOq/YU8/cXgQcagjzULNRW/Bo7FwLgQphQ81cKIf6DJ
xUq0RzQ5FafP4RVdGfAx6nunq0jITHcJkTPc9MA8seMpFXjGzwALdjQpHTI4wdExhP7rmwhoxaRKImg2k4I6uIR+qSld+IIbqqnJyrU6tuIT0owtUUO3drlx4zryJdPw
gRHnZKH7nuOp2D7SQ1hZ9k+fRJXcXA/r0d9Go+Xu7i6ih6WxcZ8uQ6L2k9gZq5Es5Fg3CslcRWCsxwMcnfzPLhfWt26e7xtK7JgVc8jStOkjPlTJc+aE7PSzruqztFxm
W4pEJhwURjpvNb0aV75pY5yf5HuhF0RKvWC9BiP0pFwK1D+KltouGncSZ3LRHlpIW03iKxJL2QQrpovhL9CD83xifVzLM35jJ1EHbliPp/1O77IR14br+YyVUlL/7fnR
j51D4xElNjYWjjvyGDGrIJ11LubQ3owhSNxZ3I55W+lZbshbc5KcF2LQznVx2YX3dhnZ3HIuCccT9ZTxmeD5TWc0dRIt1C3VXyLqYCKZAhSd66HOhArJaCLFKIr72Aws
Myf+FwN/rpY4uqy4J7cv9Aaep/1ryhdDyvSIGvfefps/XnusBxdOAV5m0MlozH3nIa+dA5BESYOVj/LmnfLFiNYrjuFA4uAy3yB3xWgP9A4gG3ogEfupxd1ZoKJBttZk
fYmY1vpQBpTvHSFIpGbaW/etSo46JNIh2FMgyDkdWK6vOBGzVRCms0f6Sl7mqGJLaYwMlnn4Fq+1WNGGpNo7LxgAEDebz2Wm+G0iH+KNpmyHVrkR+RY+S5GVSVoUp5AQ
eXrLOFUuVxe3GKiGQHSH85TPSxQ5OV3pn3j0I3adBYjR11Ayj2+WEzG+rIsIO+AR2/bKtlshAIdjfLyduhFtRhQUWfIqRlLokTuGoxi8qnYeZwTMC0/rBJXC5QKs6vNw
XbYd8pU+19Y9WJGidN7sp/VXuRioh6yW1E6SGqB9I9kPxRkMiVdrhHzfpue0WRSm2123uYmHK2mc8Y6AgcAsnM5RRr9yJu8rHAbpjIzlRSm/53cCmI5xcjK3kYi2LJwV
UB9/qOqde+mbDaqd1JX64wg3LPgoRV/dXxuq4t6hNVf+PvopMvgQekQ4xElRu4WjUOFJwZAyKwEwZu7HtI6lfIXoCcV7T+8R8i2FckZO8gm6Xrn/y2kJzQUycSVLtOj5
beOsMKn30IwMdHM2Ph4rbKGJwlDPJ2I6RZ6vRTlYsLrZu/KeLpAl9F2UYWgwjuHyXgllvTXcY9Glv/6q3VcbYcusQ0cORPw25IsZ6k8hFctCc75NpZ0lD8+ikjzwIU/b
KVkrgl+mHQLpYmwPg0ZpkLQ3A4nRPofJfVEq9Erb/23h2V1FP7SFg2nOngcuDgltp2W0PnsA4V9Sd5dO+328mgLF+cTQCI/Iakiff+3tB9iPEE+9bcXudwg7AHbsfTdw
CySh9g04ftssokFoxrc4G3YZ2dxyLgnHE/WU8Zng+U0a/8+uKO2bhFYDbBPcaphhvvb6SbdYvbah8rZSL6HChLJkSKZ64KCOTL8+pYjsFkn6QLc/UF0jv4dxYcnEsgFD
MpUjjQ60V2nXkY5MN247kdlQEMTg9MQekI8jEOr+q7GWXE4b2jIPP8igXhMLv0kR2VAQxOD0xB6QjyMQ6v6rsaIV+qP2bivj/7M4WQDvMpqXEbForzMjSmqNAS2h8lmE
nBC0CtQ5RXrX4R2gqp7v81jS54zhrOcAjw0Hlb1Y1LcMtuN3GWYlO6VA0QPpkIt4iydldj7wohBhDviqq1KbUNiUMf4exO1jSeZuVByBXWpljK9ewaYE1YBIeopCcj/O
U89LEFx9zFW7Vd3Gc9B5SqV2F6DHdvfWswl9yT7MqgI7PhXKMByD1mWP5zAXAUNelEbo2/VdQyt0vSejuamnxKan16kqYY0FGaUmYx+MoH3SC77SyJmCm6nUDYygl8Fl
y7pul/SSjKkSFppMpArJnEoFOCekFZeHYFvcr1Dn0q75iQTxWm/bMU51SUdcbXvruWKGA21NpdiCMjUqVT7osq6jnqOGVg3gN/TDlX2OQic3U1Vptlhb24CpO+NUK7/A
sUxehEhMS/LGLCtCN/KV7WTjwZHrTCzECRZLp2toLUFS/ukaj1TrgPjbXyP5Glh13yPnJn34p42I5duKUZZWrMu6bpf0koypEhaaTKQKyZyFnCZNJlVFiQA5PQKblKB9
47Ue90Y+g/h0xgK0gLZL47lihgNtTaXYgjI1KlU+6LI0pOzadPhTSD9CO9C4A0lckuuhhq4mVW1kDGh6tUBNx+jEsrowacyGp/6/k9GJnfOpeeoRbHVHBlm7hyoizMA3
yu+0QeiBLalTkNhDQR7LcdjkBSZovlqRxLySWAl0mQugb5NCX0h2/ImG4tzBlm2ATKFhubUtwAXeWmI6eC7wOXyHPixWIgAWOGUBec/OeZhG37JoTryalmDos2Z+d7EO
m9gTYeeU0JPm/IMCBezRaXnnZ63bfy8mpomRsYywmAWQ+KaeSZGuXyEAxzpRuuGVfphmSvaqgov8aJB+sQ3X/VdWs8mgMHO1AEaYGcepNGgPkfYlggKPKExota/HjIcz
0d+6ncxwP2/SN8en/135vjeudPH9serlhgwc8r+ZjzvDwhaZLSo9wlHlDop3iHwvgFKh0E2u4dtRh+pZ+S3e3vsuz5XQBj/VJuzTxOSIlhZEXIQX2dM1SfHh6iR4XR5p
xJgT0pNCgmeSk1QS4wGXgVMxyhJSAwpj8KjUw2kimH8D/WxJpu6bRrn4hDsIxZNKCqy2gTAZ/8ESgUmhl2sAPjIjL1OU/LbO2B2r4kTch1e2BLuVVekb0Xyl9Itst/a7
e7Hv6Il5kOssjJKf9XOcp3fdDwb9xCLjrsnbAJog3lU24qMHjgPU2YrwJvRG1q0iLSmtpts3zMF1qApAF06rPc3OqvbosFkAM/spQ1QrRbLRo2XR9/aWamHnqCpVT974
3vc9aqxMGeFpaENZyuJ9gJZMNnTDV+oNJU03qZ+q+m0gGjZIa4ZMliOuTd3jc8xzSjb0HH1TCjtnebO4oAM8FnTkBpTX52Q/OHkwyWCxAIqp2D8RL1+BnbMQFaoFSK2A
4p4XQ2QIrM0uIMRXD9HE2PU1vdtRhVL8t2jhUaXE3/ZTYyTerXB0su1jYcSlJ9gilP6Qb67Pxj6SFosx356NHrbjeTU9wFLKdELZIh51IdDvE2x9KdrA+nTjXyN2og9Y
UbUUtCEFEr5jEVLsj/Oiw/fmP0Y7MgrnLFkRFRnOE+l05AaU1+dkPzh5MMlgsQCK4iodqyrpkK5ghLDsNI3s7qL+8sBAYnDeYAF5dFVjshIWDpSClkZNIsHXHvru3gEl
/SDkiqkNO1sPxNsw9ela/lDhScGQMisBMGbux7SOpXzQ5lfpdZziNvOhVjrj3Ma3Xys6JsSdYbZbRp0UbTVL+O0Qw7KgWbQ6AvrnAGYyb/ClUHGa4YF0fMx+pod0kZrz
SB6jnxB7C06R0m4uR2cisgKCF3NIUvF+5TwhbR31XhZrjkBAT4K9Fu0Qt/XM+emi3mIK1aXIC1XWpQAQojC8xhrgYDkJAgXt4cQlk1/alW2LJ2V2PvCiEGEO+KqrUptQ
6by2iRKNvsR3Mgf0/cMACg2gsUZ+ctqxBxL/aTMmaosYACG4zY2L2h/IN9NrIY8uJG9z9cpvtvtgoLVnczvXtPmJBPFab9sxTnVJR1xte+uFfoGVKfBs5ERgx8BJxRct
Mm2g0d/DuowWzXfdC2XW89sQws340GaeJMAHLzfWw/XO9rxKMx1uyjBLBqQ2Ker65KVXc/wpOyelg6wbFq39dlEARl0IGTqTiVRPWzBqmztaOWrVapR9/Ig2WshrWNNK
/F7fKz9nsDQCTNzTNI5AP38j8p+UyDkmlhSueoDNYJhnHvQ8Z0kVhplr4fnbawSMbe4K8eN451NU/m/gCn/VFfVGSS72NNeWLSqIPBvh4T5kjb7owkbC60XvVJHOWzyU
IkPziNZ4ePQB/VPrKuWbZHSbgQQb2ZUnXt1YTk4A5n/kA9b/zIxD15cW9ijNhMwCPiNM1j5TB1kmTEVmEWdtOB5nBMwLT+sElcLlAqzq83Cya/dqnNjWcvNBA70X3G2g
9FcDn6YCHUMv47NsESDh8LzzFNXl2kfLvtbc6On/mIXhcs/iZXy+YiJBlzpLwkEZB0nVxy0JlfYhSVvNZo+6fnot9T9nT4z/1YQS/alwAknkgW5fFrEyA1zsFsS9xELb
OWt/aFcJU3XMQlu7Yg11TPz9ZTo9vCB9DTeueTDOU3jB0FMP+zosykyCC0XWLW24IZxzG6R8tIj1yLKly3wVn6mQsRD93GkVsUqszn74Ft9NZodwPn0yqwjmVBEej1jA
pZETpSyo4eALMFEoEHTpjyxX8zCoKxjZR42EOKNB2IZup02HJGMBTqMcCgcozr+R2lEzGrn9wmHWGC0XNNFAq45pPQOOxx1Ci+Xqh8QceriGOkeYYTotELLOsbtwm34Y
SJTJUzDhoT4DJt4vfjYriGHhgA+/DiM0DPA70xWfkUXK23LO39kRgDZn5NWOTTlpfqtjCkZyvgTZTF2HSZe8xsFOw/ifCtulZAIGTrWeZUo+iXiNjHVg4nR71olCSrYu
yogm0Sa9h4GMq195YwJtiHb/eNn8Y01W51gZlnJ8IttJYySJWlq+qXWZJR8Pwqb0bzrulEkguM8sPZbSGO4wjwGzmyL8y7f+opwcvvpad4VbJu+j8EE5xpcL0jxTuZv4
pXtR2q9zx1+qyPiGiavJqp0f31IeXI12rl5+95OeQ+oW+W9FymgZumjmQtUpnLNQWalBYcP5r6Ox0UZ0wYaydkwOLkVvBSwPjZPrhnHBJG1iTsmoKKThmcvlA5EDbmvP
zMkpd+Vd/74lO5zwiNdXOzQ/U9UL7LxwrT8AESon/HUe4Kb22cr+givvFZ7zBMLrMiw70HjXDw79vUE8PDpV9CGRdQKA6XJ+fU4VDXGy2Prdmg0z+wDvxMbhj/HswQvu
fXeIbnFBSPtXxgWhWOOLFFah3McSrjJLdz30rQTVE7NOsNsQy26JFdgjnyus/mRdcUzUUtrrV4RgaV9iZ34s36hu2eiwVUBcekKIGdtPOMD1VTH+5uM6m/REEoCTmH5T
1qclOaKrx6DG3CtnDKoSaORYqJ7VQa6RFlafG4HNBPn3c48CcDk+Zo54D8fJJYn56M4gY9ZWARBY8m/Miv6/SO0SW//ZDp71Eu0UwFqVYdS5EVlnmMZb8aw2/NQriiyZ
LULZPtAyraYGSH3OX7APeLxOHL1fdYXNW+6Vy59Q9F2YfZOScborZixGnhQSJrxzibNy7Vjv63XeUkY4y8GHjyEtpyJzxUvTubbO+dNMWvqJinw7RaFES2kiTfY1oQue
rLsCJ4obZeGMOmnz+7aU18Kj8OQiS2FFlkSpJs14bu/bmNjAg1IYfBpCGrbKiFQk9Nuqjuhy/IrhrCpHBSOoQV8rOibEnWG2W0adFG01S/jQxJBEaWr13KJ6qVqfYGbi
QFLmyM7djtjNN9r7OLqzmh1F0Dm6v1aiNpcT7IiOb8E6nU5VBhN8Y1zWRQItzeeRbXceECl6lLejzITLLSFdi42VWHnkemA9ceazOaAkQ/eyrLeDN9L8BvstK7XvvXFv
vSDoTomD5dbJPRypYr/luE+EYL7knpgePqiW0EOuGm2fBZokwhfdJQpfSPmgL+GBdOQGlNfnZD84eTDJYLEAisdBGo8oKhyrtSzcZ73RW+YzlCveq0vMQePGY8kWctn/
r9gz2rFm5xAQN9NhpxgMfM5oR2I2K1iyzuRB6WT0RF71x3GlvLNycSmJQdiSVqbU1U1l8TMeFMz+87twUhG+VGGrlsXGcZ/MwpRiKH/GlXvbmNjAg1IYfBpCGrbKiFQk
JS5kFl8ipvR8e9rNZWsGHd5OcYid6+ev7XDjlaZ2YK2Ku+t8sbYADGua3ezHvns9hiW4ssQQYBWiG2c9Olp7x+8TbH0p2sD6dONfI3aiD1hxO9d5DdKP1pgeXcW3iF6o
WTA8N86wIl2HZajD3Qahb3/sNNCWc5CAur+i9C1lPx5kCxscD/nNAZxTQ1hFB6Ey4RV5gG0ei3t5gVs7eUGIAa5XUO9BHJ5kC2kfHzI+VlmSgwHaf2C/XgXHxwdvTiMO
vzAD7RKushNFPy8xZEcfMXq2jHqek+fokHjWWPSjMrvQxI/OvcxeazATqf2OaqbT8yybqd8f9mfsY3cspq1xBIIKzEfGxjQYoa99XZaHpX/4FiQCkv5pZW8C6HR5yYB0
IS2nInPFS9O5ts7500xa+rN7NwxocI4q1P03uVhFsY0iKkqrxKOMuN+tpaJBNsOUiP7jVuaX46FY/B2KzP7BmpZMNnTDV+oNJU03qZ+q+m3+WNCKwabbQzJjx+iJHz5o
2kW67Gzwbfn/kpHIQ0o9JICmNxzirTYd7fXcs4sXVIRe3PZ8VpzFQsHkV6MewP4hcnDxWPaILTh8fM/7FSib6aTg0+G4P7aL8Qi9br6eB2FsC/L/c3ht0sddO0N2y0MR
rldQ70EcnmQLaR8fMj5WWVrUQJzqEdfc8juTcDcewh1PQfSqdu1foTt59vPxg3lYDu8ME1nPFzBvWvXSKerCGaHUyl9ktqzF3KLOGoX6Eh4ZUJXIity8A6/QxS/xwKsY
GAAhuM2Ni9ofyDfTayGPLv3vaj7+R2ADfpxibI7Ia7XGBApOSoLY3DGGcEBM9VyvFkuIuzbFohy7owv/9ddN2Fzzsg5NyAtJpOhm36VgeNRH1DPYeoX/UV9sKYxlPkn1
K8GP+E4DmH+VvhhKfWiZZUoBELkgTYRTKQljRiUfAoUeY1kqzrjGH2fcwY/D0tfEeraMep6T5+iQeNZY9KMyu9DEj869zF5rMBOp/Y5qptPzLJup3x/2Z+xjdyymrXEE
ggrMR8bGNBihr31dloelf/gWJAKS/mllbwLodHnJgHQhLacic8VL07m2zvnTTFr63v/9b2Qvum5cQ+KHA6C9mEh94lSKRPABQHkfvKJnJ+RwdwJMmZba/b7ZoNAbJJLt
pU9jG2s+QQG6k0tM+Gi0pwmMOkXoYpEqVjJ1Hm+f7+CRQ8rxnTJdQWzeSwTY0O5ISP5IZ9A78yhFoRNkBQnnSWC97zKY2QP3jtmg5o7+vAVfBdsobQlvx12GVk6yrP56
+YHgHvYE94/FKwQQ2mtpTNJDyU0GxsFi2yBUUOlmwuCY0NLYrjQKfbM6fXVP5fElnWiqPxzz5jlqFCDGCUl4rsMQaCqizvvJUSJswVy+PnqJ8q/8j3nRZpkGBik9qX3H
Dt/p2Jnotw+tvOsjV2PhPVOHZ1BvHMaR8wIn9xK2VfW7KzjUmKAyjka9giSb9tMkynABcufwcDvjK4jpFBqKuEfUM9h6hf9RX2wpjGU+SfULW77fvWcfLFLTZdIoVIqu
UN59l8csK4RAOQ+A3HFFP4CmNxzirTYd7fXcs4sXVITYfhu97vpUfr2++uJvctK5ifKv/I950WaZBgYpPal9xw7f6diZ6LcPrbzrI1dj4T363Hm5qvv+DtT/jRy/zc5I
2nl88h3fN7yp3Vsp3y0SkEPbqN0QDnow+8j5BayNcGUt6OlvimpmP03c9FFkCcPB/z/GgVVdoaGvi5l7INaUHINCHPxWW3ro8RG5qFrlYk9tdx4QKXqUt6PMhMstIV2L
GcxR5vdC2OJQB1RI6FxoNBHozJYpN+a+aNaoeQE6rouKRtkAEMylUJcwo7huOjRuMzDXCZU+VpC7FtTCgF5mjrrj4W33hSn/n2TpaNkSwm+Bplj7BNYu/ZVrmsO1eY+g
tmBlCDwI92FExkVDlKk00gfxLAvPc3zmFE4ksuAhIrl/e/yjztqURnV8GkTwvRPlkYlu/hKOsE9a2OWr5LPC4pJW12ELwYOymgEAuPZEs6TbNN+/JKn5mpCDuRztLtcf
lkw2dMNX6g0lTTepn6r6bVDT09gd1aG226tbVFjREBCPFEQW267xEJR/TSEQWjMTOm7QXvqw9nofANNbGePI/w1vdkhuprSRCZiSwoq3YXEO7wwTWc8XMG9a9dIp6sIZ
ifKv/I950WaZBgYpPal9x4okMSS2AUr31YXcUFewrNSHbEO2X0B9y7H4EnjR4k1CBCk8LgvaEZvLHm4XGMOzU+T/ohkl0SN5+FwdXSNiFiDoQLO3Sorl+HnkYiX0REv9
lTYJQ99SoTaAx1qCScrY7aFJO0DeYoPlDiZS9Yorsq1YByNQ7JxxKTl1CtbZFtaa6kp6ncrgoqvV9yseyx3W/MnKHuYsbXZwWJ5ok7RebuHDQMk8ClEpI1vDE4zOSKzs
aXisXQkbYi6jZ2ZcOQ59C7npQCE3du/nk1/NKa4qnhrR/V0GOxjSf2wFKCGDOK5oXi9DwCX5Efn4BKmi2X9BjgbZhRxQk/b115uvDVp8fYvNhvZzCqOVBx2KdGuz0tRO
h18/rZe+XKMTl+Ck8SldB7iqaRIDuuEKVcdSm224n+mQieSRPmDxdNsR9S2zblAq/l1hLstbsQGmCh7MXQO7ZmoFHXu1ZCmG3bhV3wbEcCERt3F9MrLiZrH5ZSsud7qL
WRhpwnwvXxHxhgksHVwkn1kEvnOFCdlF5bnwBZt/LilhsWwLXHAoNbyYilpKhZNluKppEgO64QpVx1Kbbbif6aqZqlinSfcSiJ+KmLr8CWzHxaBIklHEHgItPkHNu2ML
ZS9eKDWGJfKEOP3iwhVm+Jrn19oXjdW8qD11DhhdZKtvhr0TysuYj1ESI56q74VRCM/kYzhmimEguqq/NIxmVQx8HrlOafFSy62aNP0c9ArQlc64B+MFU9pxbl0XRnQw
1EZmFD40ajXoRQDlIbzO5rADwEB6rB4GIByFI6me++xWXgLvLqEgk2YnfoE2QqJ660FYLfMKg8a42H377hbK4F2BQ3hgz+JUqs23J4GHjwqwSoavkXA3OHZVG/s4ebCb
aNBKJ6iB/40Njvo4zFwPYaUzEC7Ff2Qqloob2CSqSTEgUAjyCorfbeuQ45id/HuAnmFo83c8IazQxWNbcd6dvP6+f9wl6NtQB16ZoJ37y4x0eFZqUbbTXIeYIGDppRd2
D3IJ06nQlnYSsVPNWvD2YWuITLQui88qe2A8NEMIbQUGuxVfKWEjIMt+tJKLUtk0W9ephpPD+FhPSHrAHIF1PNxRa2OXRZAt31H+07B1vDPWk5NqeOXBC9QTxYz3CZSU
dGM1O/8a0gpuuKCZYf3yKRH32UJTzNc0Kaz7n7pqBI1BO2miwnNPdKdw2YsAYFnk9Ve5GKiHrJbUTpIaoH0j2TUR6y1DNtaPTbH0Lo23oKQ75g0WoJtq4cBSqfI/arb/
zgY+b8Ry1UBsEUMF7KgmdH9BdACV2T+K1BdjHgFU51UTZMKqZ1HOmM3KrJ+L4HdD80DCUGqoDxIFiUSSSASWPMc3WHuQ/HDpT+/I+FEGz9XK5HBfR2k859hsSOAJj8vj
Ti3vJOxILZpuaa7b4E6vhiwsAFgu+ynN6Sxv+nGn4zkPBWH/FjGIcX28DHB0Vi44KqbBoYobqRLfOSsb1oXHaDiPTGN7XZR7uxbrm87EdBDfCFkdStMPCBlUZux6fSZN
Kq5vTdxpWiMagpHIEG+CcoCmNxzirTYd7fXcs4sXVIQmm5Oi+XAhKKexM+yz/b3tRjH/MO+YxPJPzCCi8KUBv6y7AieKG2XhjDpp8/u2lNf2RUbZzbZXooqU9H/jPxsJ
abGadSgmQwkNlDb2Iuw4CLRTkZtC48scT3y5SOBTyi3t1uYrn2TOsDfvGiF27MVKiaot0QAHrKgzg92tmr80UywoGt83LFHLyB4klZxdgqvB2qXeijL8BI+tsP5QWze0
O0BUPmRGPkRlEkutajL5URTDdOHo3BK2A/mSE9Ad/EsHInxiztKBdUCOE0fObmJrSjSQ/j4J67D3M2iS130ifXQ+OlzrGn+u78ATM9FGv2c6v0g9iX8yPnBxJ23aL/m5
QNAjLTJGiI4fwRdTiXS0Xy5ikYiNpSLu1/ezzjFq4+tGg0Xugm18crjVFne+LKExGuBgOQkCBe3hxCWTX9qVbYsnZXY+8KIQYQ74qqtSm1DVBq1VuWEug3d/8lyvZeMJ
WAX0aSq8jdPnfYofg3WoHSOoV01L7+igawnbk4+zTYZgxlSWq5lG2vZUg7m5CJaDe5Nsf5WX5rEpTmlrQWjF+fPGtWohsubyMY5gp5fzB4BntCppi/0uPHT9gS0fXD5F
eF70UHyd/PnkPYO3t3IoZNILvtLImYKbqdQNjKCXwWWxGUXId7FQvysB6pbmHQe/pE6YmeZIyxcwMFs9bbDg7ytywIP/LX0Agtiu7O4ItCfrjc3qBWRcbgV87mcGrZJu
YtkSFpHWmUPN9F8o8AN7KvoPMe+n2mnJ0QNRXi9IWJQ2XUTZy4bNU61F8UL+rLiBsA4T13tEiXEXaBjXgDII34GtQPQJ2wLRTcjuy4umckRgrL3bOrjUJ91cgceBjQiL
7OreLS/mhMHOcql3Zk0v0UWPGTW1qDVZ3fUtGbxb9m/K77RB6IEtqVOQ2ENBHstxV0qtsc0oR7X06bTRgur/mbelOK2Wr4KAGIiE8mASh+JdKOwO7G+90uDK6byk11xP
0gu+0siZgpup1A2MoJfBZbEZRch3sVC/KwHqluYdB7/1Rkku9jTXli0qiDwb4eE+b2c/FhwgFm76cayrLhJAPx7DSmozyUkUknixSwrj2aGBJxHb6Awuf8IUNhAWOM+a
a45AQE+CvRbtELf1zPnpopTrNA8t+HZXA0brK5a7XsrItVlA3/sRQe+PaLvyCQJzXO7hHnk/duC2aVOtdfWehmHVfQxQ0kBQxenOKGzPrhC+JG6zzXZift5o3lAtSV8x
MiMvU5T8ts7YHaviRNyHV1daHuRLua/3tZffJYtePQXcWyZzY7OHe0trPRTEPewfG2Zetz7EzdnQ+XE5H3mDN5TrNA8t+HZXA0brK5a7Xso62PxGiGCmPRubGVtJTYaQ
UOFJwZAyKwEwZu7HtI6lfKWB3+ezV3oa8h6MzPC1I55mLNVzb+wDcWnY41obtPJpbNTyQhdZ2hWpO0d+bXeYD9Hfup3McD9v0jfHp/9d+b7eGypAsnbvm4aBgFl/1SWT
7ljIPqZ3eJqV1D2w3+Vm4mTnw29GDmZcozuLu5lWZzbbqNsqP/ml/LbCb5qxET4BUTNkwM/Y/27lXxt2Iq33ih0PO8KM1PvuLY2mOQA86bykQo9u0mGhg20T8y/31s7K
kFTXiwrzVXLPni0aEIC4PM3OqvbosFkAM/spQ1QrRbJljyT6YLB6Cxbqaqs67JvPsL+l5ixmlP3W5K+q2vbiZ/U1vdtRhVL8t2jhUaXE3/bJkTx38zJquLieRZiUlINh
6YSRWej+XfI+7Mb633r81jIjL1OU/LbO2B2r4kTch1fvE2x9KdrA+nTjXyN2og9YXxL3j1TkyvfddkNO7uD1nTDvFbO3+L6gpZDZ5IjvnS8JjDpF6GKRKlYydR5vn+/g
dQZGzlnqrvykaRT8x7SiJwgKGSvYxpsqiXtoL1QWcFP1Nb3bUYVS/Ldo4VGlxN/24oya9w9tWvW4KHP8ZKPv8vDD9gT+hPD4lzesgNdTbrbhJ/GtpzphEEFLy7/0nBZ9
7xNsfSnawPp0418jdqIPWGzU8kIXWdoVqTtHfm13mA8cWdHPYxB18uMkj1Emgh2FmNDS2K40Cn2zOn11T+XxJXKHojh8FDnq9O0zTQLZSbMujnbpEEqNMe89IsafrMdU
dOQGlNfnZD84eTDJYLEAilcTdRTMEVPD/QSGv1wLnl10m4EEG9mVJ17dWE5OAOZ/QRk1UXbOlVcUdxjOQohoWhocnnT3tuiZ8o8VLBpURgSVJdnyU/Dre8ETDdm/hv+b
IY9NS5mBpbrZzCDhfZKktI+S7eUFF33ZgFTH1qwnNXSLJ2V2PvCiEGEO+KqrUptQOQvQJbABzXwBRsCMHl3989sQws340GaeJMAHLzfWw/XO9rxKMx1uyjBLBqQ2Ker6
IeIg8YZdnTAxePyaHru/zdxw11ZoB6xgIa8K+EwUWG8iMTUZoH5Ce83m3/DuwrzK/F7fKz9nsDQCTNzTNI5AP0bDs1oJVnG5qRlgoJ2bb1a0ah3bjQWDS6/45tzlep7D
UvVtURhIsJnQn98BptXoHCP46KKLdG76vlVUDOPQriDS39wPAxTAkKHH5V/BN+gf7tTtf4E3R2OzFHHxVHfEEd2cUX+kBd2DoV0AjK3UdL1EsJJD6BNHISv0xLkDCP18
lPI0k8sDounHDvEkIev1WMMl2WwB0gezOiREsn48VHpy3QQ3Eyl2fCn3sFvXPJPUG3pDuBMnb0sv4E6rkowNGqRCj27SYaGDbRPzL/fWzsocXHnxsfdqmomEYBveDvTu
UwEnK7AZiD+MRk207m+xBJ/vN8E7JB9ZcpMYc9R/775y3QQ3Eyl2fCn3sFvXPJPUtNi+zJmp/AfMpjoY8ELLfbbkdhu6xVHOQBx1EnLMK4IcXHnxsfdqmomEYBveDvTu
DCI4YzaJUgnyP5ZAQqtUe+04MWfuwcsXhho5qk6MwyzkkR2fh7tsFEruRd7sriOGC1HoHSUUKPo3T6YzWPixLuR8SgYmd/5XJ0Uk1tQPycJOpN/iInaPoj/lEtrFKZx+
lwGTxSZbB/uvgmakt4kn0dg/h1fX0Me4YNVQjttPZOaXAZPFJlsH+6+CZqS3iSfRUs7FWtjAC1ESYVdcpCAI8u8TbH0p2sD6dONfI3aiD1h1jIF1pA8C6krOFtiUTl4P
mA/1nVNH0BKbY/LPFewctKixnSrcY9feo0X9MLydn4IhLacic8VL07m2zvnTTFr63VFTlyEC55UVSmFgheMVXKQwIsYD3YZpP1purUd8LayY76i7FNqZ1plDJOzn0xXk
KWZToWAUKzEoU7qq7z0T5ypyDAfSnH2R1flpgIjDhkFnWQPfesnhDC1kb3y1s0ITKnIMB9KcfZHV+WmAiMOGQR+6rJ7Pt3a6Gzq/szqkCFvRS6GUDc8782Nxr9qGJbkV
Sa4Oc1w2yktmwEuLUdU6lJcYQURHT00uizYO1XhCtaQfuqyez7d2uhs6v7M6pAhbXys6JsSdYbZbRp0UbTVL+DpuX4a3pcXA+aGE2jdOC2+02QTVdvHB2XpEHJ7t08qr
H7qsns+3drobOr+zOqQIW/OP4rxMx2SMOcNT24JnUJWvdBDTh/4PktDrVlqWEXn5rLzPl0KNJsDoZliYcmxe7jlWVYk4Wj3I248ITXl+Y742B12IC/snA7oVQI3Nh89u
x0EajygqHKu1LNxnvdFb5m3uCvHjeOdTVP5v4Ap/1RW4/1n6FKlRVfdI000DfmeI0tRJBsJR9lc5A84p86fn3oCmNxzirTYd7fXcs4sXVISpvr2vQM8EkpWyXS3LKuv2
Gr4R8BntroPbk7kiqCzsNlV96a1t8ssGfWZex6v5PubXT4ohewVhM4bpvRq63Zq3BTHFi2lHQmkFzEb7fIy0xMftxZa2OqMcLZjS9PJtN3tVfemtbfLLBn1mXser+T7m
YRbzI2QCGEY1D+qm2loqCcmL0/Yzu/TmiE9yc9wRRv6qmapYp0n3Eoifipi6/AlsBTbrkLHwMYGEi7rgOAcdPqsbZJwybVKl/YWIiy1lHKECz4Ua8R7i34FtoCAqMeGf
m9gTYeeU0JPm/IMCBezRaa392MvEnzkc9T9bhUEWuztbNdGRdT5+qWR+7/hLWF1dEIks5L4eRsP696OBQBRhwWVnzePohoBY4aNahcoXBR0XGCnJLRgNjSSUduncWeQn
672JKnqF9K0ywnGEfJXe1TQIKm45NtwFPHNaHehu3tAhM4NjnRGkglte/9G3Y4CqULCEZ26vvOq+fadVbcJTTCP9j70699RrtmMUeior4fIBSYsgy5AAAUSjLjg2ldp9
m9gTYeeU0JPm/IMCBezRafBES3RDPXNXpFE++mJfwCYD8CxzUZ5fap0bG0O8LnW9KrQisMM79EV1kmqOMYjT7rS5angZn7pSJIRsr6bkp7ZNHgQKrd614bC3CCGVGVil
WAX0aSq8jdPnfYofg3WoHemfqRwiODpwf+joRgRZjikSkQuk2DukanquAHF6CAe3WAX0aSq8jdPnfYofg3WoHWExjc7HyKEGwiNPeBGlqzTiEj3iAcJWSeyJGc0PKR6B
X4jPGwJhI0VWzc9OiaLLtbWbKJT3Efji9Fx/97iClQPS/fgZU89NY3bQe2vmHnYivWRUKqVhFhkLTv/mXkgUTgAUhHRotNXRPHwZ2IfblKrJEDy90hBsydG01Nf3EYqa
YahCq/r0F99SYRrhyvK9UXgrRyMzrmmLjukzo+05//gJ9JdWsCXnlLGzrHJ8hwIu0Crq5hsnlOJsVJMAI3motnNyQAvlyAsz52y7FO3LfvGve4VXL4QomSBdP7zg6hRw
X4jPGwJhI0VWzc9OiaLLtf/+0cRJMwuQ1hfcMLTwuhEIt7MtgQ47GQgaCVgvSY1JMny6OPJVtssFqe4zSvn0ExwskZt9WaYeEy9uGq458mN6VNmjusnr4Vj9r15xp6OJ
6Q8BBGb8j46oeCkjVW0gqP/+0cRJMwuQ1hfcMLTwuhEVpQ6NXKi21ROlbRR/kberWAX0aSq8jdPnfYofg3WoHbtVSLu1PPATNfivLHqck7w6mbDONG1/NjswJkNwITTG
yu+0QeiBLalTkNhDQR7LcbyzwU4GQEBkMt3M5hFbrKjdFs/RuAxqjCFD7sSwdLNu+J9h+KovGBMCYQa/Mj5O95QTlsQojoA0N8+GkncyK3YHdqZqtqxaQ8nVKdJdvQCU
fphmSvaqgov8aJB+sQ3X/Wzkc6+eh8GdIlm96njmtfl9U9rgTk1Q16CQ3WEIhWTDOz4VyjAcg9Zlj+cwFwFDXvpclbNW8nKFoYSzDRdgXrbvtcHYUKpXp+rzYYxS5KGu
dA67pSE4aiz9sn3yDWrgH6Io6z/DAs3VtaN9ZVXI+iVayQ4qXvYICukxcNFd258HY0NRxUENtN+zfT6XPmFPORyMr/rMOrct9EkrwhWenz1ifkkA8Ao+sbZvntLVJsKv
uu9bgvwv8ZLc0NjXWEfDDBwskZt9WaYeEy9uGq458mNn5iCzDf6WS03MBocytX9UqVu6MnaBCMysuW8+bF32tP/+0cRJMwuQ1hfcMLTwuhHm5QdVPr/XIfGZeYP63GuA
EIks5L4eRsP696OBQBRhwbtVSLu1PPATNfivLHqck7wPbHyOAf2TldstJsXcYBiExJgT0pNCgmeSk1QS4wGXgUkP8TpzzQ52HDRzOcBWFp7H8m7QwCRf8+XfYAq7Nc2X
lbd9eWkKHkLUuzGOzBgOG2zkc6+eh8GdIlm96njmtflfu9j5US5/fWMkkaCP9xYUlSXZ8lPw63vBEw3Zv4b/m6Io6z/DAs3VtaN9ZVXI+iWVySLZ1pJNJAqwiBqbf24k
LmKRiI2lIu7X97POMWrj687EO8/g9uwsqIMhrBIGwi5HcBxv9kzzAGzz2DaA7v/Ba45AQE+CvRbtELf1zPnpolLvzXILZF6ZBj4xpTeZd7Sl0VvdBTXNh35mhVwSmpx4
47Ue90Y+g/h0xgK0gLZL45so2n4xO7x51F11DJSw4XqLv0DXTm7nHoUN6iiCY8WtU5mwg72j/oTeW5zYyDUkVpso2n4xO7x51F11DJSw4XresqQeWApN5Y5y3PN6TpUZ
tvVpGoJWHnRYEPOGUh6p5c7EO8/g9uwsqIMhrBIGwi6kj7QSJ+cYT8iTeC/rcgLEUU7DKFPHlwM5NcXgy1ELlpso2n4xO7x51F11DJSw4XoNHbsLSRfUi5XD6Z48kp3b
ofu16oqgy0HScAQD9SLEa1LvzXILZF6ZBj4xpTeZd7Rdax9/rui8Hi1KcsJEuFKNHtsxIBVIgs4lmzBDcgZK2VLvzXILZF6ZBj4xpTeZd7TXzV2JgtTyuKt1oK8tAVUf
+YkE8Vpv2zFOdUlHXG1765so2n4xO7x51F11DJSw4XoWANpyweTELwMrclE510QZHvEwJCHh77CYNr7vwcFbApso2n4xO7x51F11DJSw4XoRwZQVFvJr1erL9ezYf7Yv
5dWIQeFu4DCLJTVajfUwu4PHBXo0Bws0nQo0Cu8Lza+6Uk8v/zUdnh8mPOnpzqCAbUZEUMpCpuoE78yr4FEt5Jso2n4xO7x51F11DJSw4Xq8RzMVr2orjFn/j21Y53V1
a45AQE+CvRbtELf1zPnpopso2n4xO7x51F11DJSw4Xr+3Vw39MqJtWrtekfaar/6Oz4VyjAcg9Zlj+cwFwFDXoPHBXo0Bws0nQo0Cu8Lza/N7lFin0pQdmlwobUxuvb2
lSXZ8lPw63vBEw3Zv4b/m5so2n4xO7x51F11DJSw4XpK+9FjLc+usCPW9EhhurT7Gr69BUVQlXIVeJaZZKOqvnALloFM/swh6ne/8rkAEtp/I/KflMg5JpYUrnqAzWCY
z2qXRnSx12BqDmkkee9QWnzhubEuiOa7CJ5wDwQF7gvN19is/npKKV65Y7oT5mrHIvd5pe7CpMJl9VPH3AdYjRuytIWc6oVaWvfP6br1g1G+JG6zzXZift5o3lAtSV8x
//7RxEkzC5DWF9wwtPC6ETdMkeXKMLeAKQOua9Z75fZYBfRpKryN0+d9ih+DdagdZWfN4+iGgFjho1qFyhcFHa0mGtFGJXE8e8glHmxHzUZQ4UnBkDIrATBm7se0jqV8
MJ4FAZzeYsv4dDFgwFrDsniqvOZLZFTDZ48tD/6GFk6rG/1KimxolJx4MB89EJ2XPNCVzcWO8rRzPyQISqAE5VIGASDXJ+j/e7SpF6VUXtPK4Gz8FFMSXpZIKQAOGQzT
OQn+z27saTsf5/vBGJysxoPHBXo0Bws0nQo0Cu8Lza+ZsuDelh4ye/LvUT1wCknCa45AQE+CvRbtELf1zPnpopso2n4xO7x51F11DJSw4XpQ8N8FFB7e2ASKv2lT46Ro
Lrr5p5sPBZTsqoY+RQ8v+ZQS8063fI7C/ueRb/zhZSYdlvk3HWcIXs7f3fPU8v5pWn3naEeVXuTMadcanOpUc7Ut5Y3Rtvx7j3T1s2+1zJXpDwEEZvyPjqh4KSNVbSCo
tQhdK2JnrHYTPgMm3uzNpVlTq9qbNWpiaPsK7Nt6BQRQ4UnBkDIrATBm7se0jqV8rf3Yy8SfORz1P1uFQRa7O2kMkZNtRqLqeNHJgMj5ZSXe9z1qrEwZ4WloQ1nK4n2A
GzV2A4TGwgI3XATqn+uZrKpmJPGceAeuncp9a3gxbfdrjkBAT4K9Fu0Qt/XM+emiGGQHJrGpC9yRZNsQGzRuLlObH6yLLgULvr2D9+ptfVDdn61KE6lRri0QqaV6/H+8
QigO54lGH06KATX1Sgt1Fx+R4H/oikmKchTemGSzYDWBfhlLJwQB/JSp3lQfz/5dUHLfOBqdG9QLO9Ya+iK5q8bqxvpb66XJKdKn8TQEjC3+copfxFWRGNiQiQdTvPx8
4KU8pRiQYkY29hI3F7dMlLqIOBRwkE27a93xbVamnCHdTwnSf2ocI2HNEhWWutzS/+2XQ4i1rxW3xSnaVXupUNOQ8YjoAko5/SSDFCnh4Ok2/8G4SJVd/UsKatWyD/KD
GKMq7bw6cyYqBSLP3fllRBA1ZQEX1kTlZO9tiHXVpbpQ4UnBkDIrATBm7se0jqV8GJCKhVWPqWAsY4KpVwW9qG2X/Y2/6SwkmuCmwqbnDr7LTQKawyhWTq0qzQZ12mUb
w/W6SBrSGGb4M4TJ2SnbwhWp8Logo3lVQP2nJWLnQ+EcWdHPYxB18uMkj1Emgh2Fm45pDpHNx6cdEvB3UxpBMDdd3pJaJs0B8IB0E3BrzOSBfhlLJwQB/JSp3lQfz/5d
1Ght58T1Eyakwb01Q1+RxmuOQEBPgr0W7RC39cz56aJMlgQFDS6ZHUBK9BZUNDM3E9+4BAOMlIlNuG1q3DJWkM3OqvbosFkAM/spQ1QrRbIE6d9w20HgOWHZF4EYKRR7
ZI2+6MJGwutF71SRzls8lD/v1K1HanNjYYKo4jnZGxLG7xWBEWDXZNQFTaJZA6/pFt+XmRlL11qhV4D7fNe+jKOvUGVhZMGlmBYgnKRs2qV1L4jdmutXmpoS0KWfLRN4
hRzDBQbFo50WM5tCM1DxJro+Ynm0+3sGvpfShMGCxCF8hz4sViIAFjhlAXnPznmYm7UVtGXgtsZJOEZBKCo/hvifYfiqLxgTAmEGvzI+Tvfyav7Lk6e3IFACMt14mh4u
KbVwFv7lmIE483NxjEeS0Vzu4R55P3bgtmlTrXX1nobVvH72UR7D40czmPiLSV3iyu+0QeiBLalTkNhDQR7LcQfG6m5gv6+xv/+xmiIt8C9ayQ4qXvYICukxcNFd258H
N+6L+kQ6csLvVW6r/ooN2iK6SE7OHmr0x6GCsHaazRBiLeyb8ViQs4vr4f19RSjD+J9h+KovGBMCYQa/Mj5O99ns3NooWFPU6E7h7aeMhlsptXAW/uWYgTjzc3GMR5LR
XO7hHnk/duC2aVOtdfWehryCZqw3/fMC5mzOsMf6g5rK77RB6IEtqVOQ2ENBHstxOK5e6HVvBbHLmtvLx0unWUcmkr/qfrp/FKaoUcVT0v+UJ1Ia9WeBfVq7EAYcDVfA
uoSsBipgRnaz3Gu1CZPTDTfui/pEOnLC71Vuq/6KDdpN3PqA9KUmDfjTHs1cMCPERQbuEhtD/hz6kjpTD+B3xHyHPixWIgAWOGUBec/OeZhwugNNveV64sPweHIK2ZHu
+J9h+KovGBMCYQa/Mj5O99mJHxwYL95xIqnL7VIOKIxYBfRpKryN0+d9ih+Ddagdy+/KBcRvy6e+qn/l5K8lCgRqSZh18P0Ma9yzDYmA5gDMB+9cadiOnkTQ0lTocvF6
0FivrvCLnGLHeDBtfnY2MHSkRXWW5EN/fh9WHrVOHkWQ3U9q3FAufoBEPwYYR/v10hw85AdyaxwRVUL0/kXX+sqIJtEmvYeBjKtfeWMCbYj7zO8wpNZ0sCokNAzPLYPw
LyAFnLQrQDhbvS3+nJra0gYizLDg+LMiXH0jd3Idj2IGBBwjXLt3NHixMztKf1vhXUFvmT7r0ptzNDJyE6YxpDEZbFJXs0QuBFtOmraCeW6ShFEPum5NWjpCgqaDqsAB
rwWHOciDPtnhAH3ob0p6dPVQkfyCyzrIrzvJJweBX7U21edd5XN/3hBGKeSz/jQR9+GuRMfhV2pb5nqwsPi6GN7YN+iWSI0zfA+1UPUf1bKCepKn2NgEZy7mYul1Oe5g
gwK7tNWxHrdLW3NDSNqCGt7YN+iWSI0zfA+1UPUf1bKCepKn2NgEZy7mYul1Oe5gp7To3mE57UsS/+RBftvPJt7YN+iWSI0zfA+1UPUf1bKCepKn2NgEZy7mYul1Oe5g
85pzSd4//riP+vBfH3zcUy09OOChCvTVohUb6mU5cMdZAQsW/mfx/ZM248LaiUvIjXZl7tAbXOkUgAfAtQTFveD5JUMUbKwmnEBIBoIW29lSj6m89qTLSKdC7r+X7ex/
XhGf7mikKVef0telrq/m2n+kCglz3xLhE9yxpeI4zEP1B3Q0BPXEHlFsn2zFbSStq3J1SjMH1k4FLkVcmJSM3Z50gqo/dpuZOOwI6c1IvIdYGSdKexwxz4j99Wn3RD+E
HQ5w1eFb0JYTrKrbUeNY5j44HmBoO+Q+jYGIEy2FlsIFOiEI6xbXtJYrSb1j7dm1zQJwZqgzNmUmTaIIYqV1O1kBCxb+Z/H9kzbjwtqJS8iPmU75KLAehQ9j4sNOEh7s
M2lbwi7q6ZAxuOkVWp1N+B94qQ4L7qxJfqS7JzahDQenqVHzvrJv5B/sgErAnBd4YJvfskaxJtOh3oEz4FCQL8bfcwiuz5bPOHXbYL7JlXEI4/CB9Kx/KQ2qjle9u7oa
DNm7D25de3AsJR/ZOicxqmyeMO04ZzJCIES3tO1izaxJYySJWlq+qXWZJR8Pwqb0rggwLrGV2pVqBHbWejMPZKPKcDvpeeF/LO/+ofJp/xfe2DfolkiNM3wPtVD1H9Wy
gnqSp9jYBGcu5mLpdTnuYKRTthvASuvEARZhl1AmVvnP7QrSJhQxDNBQupkyF9+BG3a+UcOJ8G46xR9nV/juzZJ1wJ8sTHsg/qtgo3hp+e9sN0U4JAvR//t8wr4q95qp
/o5/b/kR40fauObkKvq63pDdT2rcUC5+gEQ/BhhH+/XIddMVpKuhBU6ATsLr/46Cfv3Gij/pC7X3nzbuBUF/7yTgMk4XjNz7CIfPz+6cVSHKiCbRJr2HgYyrX3ljAm2I
qT4fCpsUiI125SFiSA0PNq3F75sspHOCwJ64J6v6T1IFK5rgym9oi2C7DujpkuvKN1MxHoGEmWcZEI2uxQJ4Fx94qQ4L7qxJfqS7JzahDQfpc7X9imkMsaJypTrb3os7
qf3bRtR41YSzfsRhNOO3d0pgL42hInILVL6deCItikmCepKn2NgEZy7mYul1Oe5g+PB8w2FAcSpQL6H5xGQkTFhpZ7LkOMd+g7VaSJ+YvxhC2SZ8RS0ftOftsC5mfZf7
BiRnUo4xcxjROfQtP1jjfMW+v893AwXKS2So7mgMfces1hAQxZxtKLBZ7uYO7stYSDvlh7QcoTNYSZsHnlUPduQ6xhqaSV8NcGaJyuRT7IPGuqUNEUMzhV6SQAWg+CF1
gpZBSzNKBNXcraWGJROdJxTja6+AQstXiFdZUst6IydemUCObMXSpWQIMqKmJN4ESiGdAIboKY9SXPzUKSG4Wxto1TruR4eZ1tECV23cD25/8FbGTmyEko9NwfApVa0/
RMe0g7shdEuSAHNcBohXCak+HwqbFIiNduUhYkgNDzatxe+bLKRzgsCeuCer+k9S3NQK6rmU1MZeJ9AKu0dgWZJ1XxYpJ4CBzJILILhMHsfRykurN0v+m20WOq56XDJC
fv3Gij/pC7X3nzbuBUF/76F170t8MQz+EmGyPvkFFcapBKH2C9lbfAk/matsO1NEjojpSxUDID/t1BMe5UXdqMa6pQ0RQzOFXpJABaD4IXWClkFLM0oE1dytpYYlE50n
FB+OiPSYyE55etxBaeNGbApS60pkUcR+99KnH7K3C0eqr0ZTEBIJNM6Y/crWOEzRbztmR78bGJkkrUx+KGBxjyAO+1hXMbvHC0qlIv4w2KKWR+JWi6+ySV+A7JH99vIe
gnqSp9jYBGcu5mLpdTnuYPjwfMNhQHEqUC+h+cRkJExqkRqV8SR32fpj/as3J0R+kN1PatxQLn6ARD8GGEf79ch10xWkq6EFToBOwuv/joJ+/caKP+kLtfefNu4FQX/v
Avrs1jiUib9Wmq7zpi7SFvbeshtcbJO9GascshhESO+pw/0g9BTpjxtq3fdVjTx44buRwVhLdfLrgVnZx9I2k62Jsefd6Qwy3BTLGnHfQcpeEZ/uaKQpV5/S16Wur+ba
B6wyaP0o5WPZ25IoU+tE9rN7obktOWkg/pzBD0cg49UNg2ydJdNhjlLcGNXUFOTlfRwA4CIowIbvCTPm7QyoWD6N0bCtm3dBOYx0FY/yu9wxIaNyNYfe8ZzGvK/qK3/D
JUEtjzQRd7wSfboWHP/B2KdNG2tI7fwxIiuSthHusS/bBlD3tDYWCrIlMmwZUq6qH3ipDgvurEl+pLsnNqENB99VD94fkvjyTq5So3V+89vdN18aGfe/vAcCGj6yYBIM
UH8hFfbTRe9Hg48m2/5XwQYkZ1KOMXMY0Tn0LT9Y43zFvr/PdwMFyktkqO5oDH3HdOwG7N0LWl9CQv9bVzOqI38XC50MpcqcWZ0S5gPd4bCedIKqP3abmTjsCOnNSLyH
9+gpKgS1cBvPR1JCo3PuAETb0PckcayTEhQPYxa4EfD5cLARmjoPf8KXhOSKYTBzfFG3YvvZYhrNMZ6NsABjAeG7kcFYS3Xy64FZ2cfSNpN6HEmHbp4bSK78DsATTTTA
lxgvC4Amm9cQz4dvxVtCGc/tCtImFDEM0FC6mTIX34FZAQsW/mfx/ZM248LaiUvIhLFEsuSi05pIZzxqztlf8Ruw6b22lVHPXwJOMPSyVX9C2SZ8RS0ftOftsC5mfZf7
BiRnUo4xcxjROfQtP1jjfMW+v893AwXKS2So7mgMfcf6VrJFPClCtHU/toEVRssKCOPwgfSsfykNqo5Xvbu6GgzZuw9uXXtwLCUf2TonMao8Vd1Vu3EV6klk/rqD+dUq
ooelsXGfLkOi9pPYGauRLLZ1wTSsICUeTq+2WvKbUdR18CQZSHj3HBUH/hSRrhTNMSGjcjWH3vGcxryv6it/wyVBLY80EXe8En26Fhz/wdha6aUKufAb0zzGn4rntwbo
n/hpH2IiGpTMsGN8lhPt71kBCxb+Z/H9kzbjwtqJS8iEsUSy5KLTmkhnPGrO2V/xwfBBEeWgevRm5av2+damaa2WPl3UpB+JWOqJkkljU1euCDAusZXalWoEdtZ6Mw9k
6L+E7lZtFVHIJdIvKyg2Cp/VviaziMebYOWC52xAWw1n2ZVPtJVGiEI0K7PCiSrCyjPSRhvsH2/7PvdLVgV2csqIJtEmvYeBjKtfeWMCbYipPh8KmxSIjXblIWJIDQ82
rcXvmyykc4LAnrgnq/pPUuPCy8CK3u76S5FpvNqFSePALCUnkOIcNL1rUQFp3eGLCuNSGggwxVyUPo9RUQBHK2MSeq6kh/6a0MiBjU7eFkkxIaNyNYfe8ZzGvK/qK3/D
McSWsKWAChUzquZEtP3a1/kfXy+/CpWDcgpXmK+zeKR3KxmAGr9BoVcuPk8HgRDB3eG/YpXyuVJkUi+vhyouiu8fI7rwkHYAlc9S/F1McsA8Vd1Vu3EV6klk/rqD+dUq
qcqXXbDf9GRZdsbYfOslIE17uyQNL5DqRuV3Wp+ve05/sE6BNN+3Ems5VGt1qP2AR2xPEdIx7xRpEQD2z8jxgc/0maE1Gk5bIM5MPOWOSiLMB+9cadiOnkTQ0lTocvF6
UfxObbliAFEGzmkR0kXwTgW7OQ93GCpxKsYB+PPnstvLtxKF8BX8MTWfIP/0yon3dtjJRmiIeBVC5578IXjZdChUcgoxtL5qmxVnrMJ7+6ZVdIZ6YAWW+eJSVFvyvMoR
i5sEJDsjSGyszwCXMa1kLtXJvF0jVKdLjFIfezjK2L4qQdNgtnd4VWBHoVyrxvysgXHzJ0vhCIY2L1v8epdSDQTW6n04JieJhfeOesh8Hwr+fUVLe5hL+IYHzPnwTPG4
BPhD7gRp3Vity+ehrhQss30cAOAiKMCG7wkz5u0MqFjP8xGdbXzAZgJ3C6IeZXDhXlJJHgXu3nbjsIhCQtevNV4Rn+5opClXn9LXpa6v5toE2SBjoLAO0UtN2Mk/bqWE
t2X2bI/12l6Xb2UCIWdAZ3m4q2SHPiHMZfBUKInVcFgE2SBjoLAO0UtN2Mk/bqWEA6jWyvz8ekcpqwhUHJhAfkljJIlaWr6pdZklHw/CpvSikTVKTJI1WRv0dbWwnLb9
pgeI0frX4Of1tvxaB6Fmkyt4yzJRwMwbtPp+vPYF5BH48c7Dt7hVh/xmGb6ZkmBKMGVvSxOTV0mLVRH+v8DWyNJMZ45uzt8r0f/MToicFDlZ3BExjngs2MIk7MHeXB7Y
YrYBYJNIoFZ/19GO7/0QYtba4Pa4NYH+wm5p1i+Tj/o4GBIuA+CKAb6B1H86F9TeFB+OiPSYyE55etxBaeNGbCMTUsuHPZIoa8u5nYA6dinT6ZJKYHskXjmKlELUxrHn
tnXBNKwgJR5Or7Za8ptR1GctMZUltvV45qVnE5Y5Hsk7X2XSy3mfgskI8jTND5SX7AYBgWZTv0w88pn+3PicZVLPVvtupEaIAYpwPbgqI/3xtAHe3wH1gi28sBhXJ/sV
OVsN5v6pP17OQWUf7SJNEG+/JrZguQlNWjAxQj1AHS6GGJrdhV+rSsyjwxS2ocisi5sEJDsjSGyszwCXMa1kLrQ0N5MZoPT3L5ZpEc/eFNKE3gtIYGDNgDcBqq8eNgMj
3h6F+/Kx3+rXKoGLo2115viKkp6cX9upuTj60tlNg1vE0AMscUyBA6tyq6FbdyNpOEOspsrUYKuqco4yRpah0gWmsXj2ah0jEAWK/qPR0lXmjYZGTPpx5fHkDH12aeTG
rKB3BhrifOOJCen9A1+VJrqrgu7gFnA8p1pudqBB180NqhPwD9RVy26NTbrj5fBFrKB3BhrifOOJCen9A1+VJmjJnC2ZcqDo9Skghb1PLQam8Q0zWoMhw0KIIPISa/45
2MmhsnNAswMAwHMvN7xnlhSHpRaErirurfF1FNRgdLp+6NLQUFfar9A3HyGbRkeiXxTyWFdx/vN1dPovi3M8YGqEuYykqTsrgwmmeO5vcDiRbbIy+BypJuhmaqcoXReT
X4RQscDfrERbv7VGPOSaZzWGrRssoCB1nVcRteud/OF0ecFsytFfT5AGNCEJWV5prNZyvWO4V//x/oYGun0l/kyTto6znwCQBLvDgPsDSXME2SBjoLAO0UtN2Mk/bqWE
x/gQQ3pq0wcpSAlYYJixiUljJIlaWr6pdZklHw/CpvQ4Q6ymytRgq6pyjjJGlqHSjTzsfYt+G2EtkSKdO3dkJcJ4aVU78MKCa/37RhMQ4hMUHA9aLezjViBp0xdmJs6i
hnK56BRUgeX46foVuyM+cN7YN+iWSI0zfA+1UPUf1bIscjoNBMu1CLtqI8qHDyz5HmcEzAtP6wSVwuUCrOrzcIsCv/DBYlaHOJQLOWWUFWEk+xOpR10+rMybAicjUDZS
s3uhuS05aSD+nMEPRyDj1cWGSAqgRrQelVZzrI6erO4K41IaCDDFXJQ+j1FRAEcr2xvaQ47JOsOhci8Ow3+llTEho3I1h97xnMa8r+orf8MxxJawpYAKFTOq5kS0/drX
VDG6VM9urcNjt8zlDJyeEC09OOChCvTVohUb6mU5cMdZAQsW/mfx/ZM248LaiUvIhLFEsuSi05pIZzxqztlf8Y5V5UQ4tP+KBUx/shTz7tQEVdKVch5YWxhoy8dyuHDt
1iLUI8jgDTmXmQ3g4KL12OG7kcFYS3Xy64FZ2cfSNpOiDFeTGUmz2p2f9KodTz4Y01p7wy6h+2IuEeIx4RN8F0LZJnxFLR+05+2wLmZ9l/sGJGdSjjFzGNE59C0/WON8
xb6/z3cDBcpLZKjuaAx9xxIsH+XjnyPGSgFEm7/bs2+6q4Lu4BZwPKdabnagQdfNDaoT8A/UVctujU264+XwRak+HwqbFIiNduUhYkgNDzatxe+bLKRzgsCeuCer+k9S
FdgZUOlDOkKFY0gROzrVxSokUTyqZ2mdegnUq8OLVEqMPZbYCTsmb7i3kW+D1n/R4buRwVhLdfLrgVnZx9I2k6IMV5MZSbPanZ/0qh1PPhjuMafyjgLy9k3WohSpfv3f
3rdgMwHcs5xHKxXHDvdw0NHKS6s3S/6bbRY6rnpcMkJ+/caKP+kLtfefNu4FQX/v9x74S6WiDokmUgbFKtopLzBlb0sTk1dJi1UR/r/A1sjSTGeObs7fK9H/zE6InBQ5
gnqSp9jYBGcu5mLpdTnuYPjwfMNhQHEqUC+h+cRkJEyfDEY0uJ6ivSNkcxiiJZYHFeHxVpPSf5PH41cKfri416040h5ouG8/9bxKZBSiRBJKIZ0Ahugpj1Jc/NQpIbhb
XZFSQgg2YhncbxqeMmnrMOMY8szjD05s0mWan8C0QqoI4/CB9Kx/KQ2qjle9u7oaDNm7D25de3AsJR/ZOicxqjxV3VW7cRXqSWT+uoP51SqpypddsN/0ZFl2xth86yUg
1D3ykz9mrBRmRcH7cLSu1x0OcNXhW9CWE6yq21HjWOY+OB5gaDvkPo2BiBMthZbCbU9Ub95AzUy2zeLfcaiG2upnm+7tWZt/WupI2zb/WfPrI/Z0xYgFH/C9SJR6H/t9
pfleYEHmnBrQz5xTB3yU+B94qQ4L7qxJfqS7JzahDQfEwojykNOwdMABhr1HLtqbOeMNQ13uVwgVEpHKmggJcQInllDQ/LeNQQC9W9SrcOVskeNOkxKL28ryPlYQxDDH
rZY+XdSkH4lY6omSSWNTV64IMC6xldqVagR21nozD2Tov4TuVm0VUcgl0i8rKDYKn9W+JrOIx5tg5YLnbEBbDQVjvjSpVkSlWtIGLmYbnb5HbE8R0jHvFGkRAPbPyPGB
BiRnUo4xcxjROfQtP1jjfMW+v893AwXKS2So7mgMfcf7ZigYx3D/J/uOoduvkkLOsncpP6DOH0G8i/7wsLkgwU+KPsnBYzS2ovnuXxWVg88+OB5gaDvkPo2BiBMthZbC
bU9Ub95AzUy2zeLfcaiG2hxT5WFtOBA5wmMVie4VjMelrPScVxFAYDUIsn8iFNbUR2xPEdIx7xRpEQD2z8jxgQYkZ1KOMXMY0Tn0LT9Y43zFvr/PdwMFyktkqO5oDH3H
+2YoGMdw/yf7jqHbr5JCzopsAsrlIEic3TXVp9ZnAcpVPZfRK62p1cM2QSUoF53Nafcf01YpHTUfhdSkhBxEmCT7E6lHXT6szJsCJyNQNlKze6G5LTlpIP6cwQ9HIOPV
xYZICqBGtB6VVnOsjp6s7ndE48XHt7GBrIzJf1GPtsAtGw0PCF1cAUm1C+9L4u3KvbWNJY6eTH4cqDRKSZ2uQGMSeq6kh/6a0MiBjU7eFkkxIaNyNYfe8ZzGvK/qK3/D
McSWsKWAChUzquZEtP3a1/kfXy+/CpWDcgpXmK+zeKQf6xWa8wqk0AR+esHtnsIZwvo9j1w0NKW3ayatzWLkCcuhB1z+K7F4X5y5WUUz+QvGuqUNEUMzhV6SQAWg+CF1
9l+rTswCk8J8vFuGT8lLhzd/Xh8Ufzr/DZwvjxoNiEbDQJOtGbsRnX+5a3hR3YuaiYA3mjgttDnv99OUpr929hLOnup52fOeAjXg7myxy0+qr0ZTEBIJNM6Y/crWOEzR
Kxzrje/F5wU1J9G1vZvdXyvbkWAdTBqT9jnZgr+cJViZdBno9IR1q5aM2xYYs3rLqjBlYBfZH6CM4IMAWCDpacJ4aVU78MKCa/37RhMQ4hM+OB5gaDvkPo2BiBMthZbC
bU9Ub95AzUy2zeLfcaiG2hxT5WFtOBA5wmMVie4VjMfvmENKZo2HUYjn0uzoJFTg+j/NiNS0Z0AmKGf6UrQuPClIkOjXuZK0DFFus5b2QZOf+GkfYiIalMywY3yWE+3v
WQELFv5n8f2TNuPC2olLyISxRLLkotOaSGc8as7ZX/HS9DclKqpj0/hxCj1or69pW5XAmUoey8ZR15z3OAnz4y90M/V9SD49Jm1GvE1wBiq254NMbTZ5Xf3UhC45u4+p
zF+bhteOBkyb+EE/DwL4YkohnQCG6CmPUlz81CkhuFtdkVJCCDZiGdxvGp4yaeswEsQZI1smfWMLNvbttwQXB1+g+ahR9MomsztQdwoKfHvqMzpgsiGwRi/aiuY6xNIp
xLwhJXN1ZtT6cOzFD87K7tsb2kOOyTrDoXIvDsN/pZUxIaNyNYfe8ZzGvK/qK3/DMcSWsKWAChUzquZEtP3a1/kfXy+/CpWDcgpXmK+zeKQf6xWa8wqk0AR+esHtnsIZ
ZQUNydii1ARvILmT1ebO7LpGPjWm9Td21xrd4STsflqBdJN2EA0AjFxAGDkQjfpZxrqlDRFDM4VekkAFoPghdfZfq07MApPCfLxbhk/JS4c3f14fFH86/w2cL48aDYhG
w0CTrRm7EZ1/uWt4Ud2LmilclqekI8wW3qkvObf1hTsqQdNgtnd4VWBHoVyrxvysgKyeGpX+/UJSxYqmclei7tqKXbwT337CD9b+4rbItHwK41IaCDDFXJQ+j1FRAEcr
A94Zyqf9REzG3RXdUDRDRxXadCrg12qe30rKQeaQEgl38P4fd6BXNxcLkb+4Gl6F41FnfCeZkFJmaJwalVa5hBpJaNdLlbqcDCsb7yLmECNVFOFuvZEs1rY5Iir/yI7U
JWqbhbiJQgB/qil0YMty1HXwIIj34TbQfcM3X8/k502Fojm84KtKFCa7mhMeosRJK66wtO84fnWgKZggpMzpbW56aA9lNb6i7LrJ5VJcMstagDfPXq+JsDPQKRhH9WyM
QJycXyaECaoVElPm4eMTfqlKQFjYl7qXGbSBCXmVGv25jnP9SIdSrCwe+Y6uV6lEDBz5Nr/AeyKk5FM+5ulvc/0DHNe8CgAADUqIIZtuE0rCeGlVO/DCgmv9+0YTEOIT
mnT7ks01CExe8gDk4koafwVtkgQSP+MLt/nE8ufbJbbe2DfolkiNM3wPtVD1H9WyA1UdnG9Q4Sl8nnHOS5G76pNl2oIOSOD+xFBRkhqDPfmLkil0UJwP4VVNvOw1v37Z
MFKSLIQQL/2TI3aRLBlKacJ4aVU78MKCa/37RhMQ4hN4UrsuTYuzK2V/z6ADlk/9kN1PatxQLn6ARD8GGEf79ZCKmSk37yeBiOtQEgs4saERpLOZO8/5I4tMXhiHb3U/
LCYYfiSNf5qbH0HGPaXe47N7obktOWkg/pzBD0cg49UNg2ydJdNhjlLcGNXUFOTl1/nLfe7GmLQqVF4SdsAoF48ulOhCEuiafI0XOkb2KQThu5HBWEt18uuBWdnH0jaT
ogxXkxlJs9qdn/SqHU8+GLZH2NSyZf9bpQIFbKpYjYkK0hDruhL4VzWquFL1GbXm2kaS4KYyLN0MGkjgsq43LFkBCxb+Z/H9kzbjwtqJS8iEsUSy5KLTmkhnPGrO2V/x
0vQ3JSqqY9P4cQo9aK+vaVuVwJlKHsvGUdec9zgJ8+MvdDP1fUg+PSZtRrxNcAYqRvElZ/nNEvin299h7hFVrBR4YSI26WYsdfqk897sE+CeCpNZccTnOF6soZI82rsJ
Gxl57raIGU4VFjn4HiYWbXh9d9Z2Ypn+WHfHMyuaAV7k1B7uR+M6RBtW3ImmghHR3MdtpeBHfo3NG/VRFzD8lbJ5XcFYT07H3XqQ+DOz0UnZXHKHmTFCVAz2skLnLZ3Q
o4zufsiewE83qecRKB0IQo6AXnezkQxRfaPf5W4eA/r3sYq8670mT8XihyNiMze8vQzBqTMoWh/E8qU01s6QGMPMURu4d6qRcP6Z0dNv61vVybxdI1SnS4xSH3s4yti+
yogm0Sa9h4GMq195YwJtiCmwFpr7r3fIpVdYnA1fXcvOKXkymeIWk1439kH/fHbZRAtawKFbnELU3aPyIFnrGVkBCxb+Z/H9kzbjwtqJS8jGv8jyfHPIiLSdovnsBzVm
ia9fmNFgGjI/5LT99C91GmQTSgKPN2Pbyb+8iWDdTcZq6RbqOq9W56mAGSiv1b8sOBgSLgPgigG+gdR/OhfU3urOex83Cf2TC7EyD9zI4+ApsBaa+693yKVXWJwNX13L
ZBNKAo83Y9vJv7yJYN1NxtvO6Z6RqaBtSwQ7p/bpySE4GBIuA+CKAb6B1H86F9Te5n3MAXeRABCtO5IXt9wC+ymwFpr7r3fIpVdYnA1fXctkE0oCjzdj28m/vIlg3U3G
9+XUCxfGjUIlDC4Sy094xjgYEi4D4IoBvoHUfzoX1N5/qIDNIkNHL+CH16S3wPscKbAWmvuvd8ilV1icDV9dy2QTSgKPN2Pbyb+8iWDdTcY/d77q3/9EHz1jgr0LYHg8
OBgSLgPgigG+gdR/OhfU3kgDEI/1njLw+y/b9uyHzaYpsBaa+693yKVXWJwNX13LZBNKAo83Y9vJv7yJYN1NxvjbPYPEvgBp0hlaCd+IDyQ4GBIuA+CKAb6B1H86F9Te
x7Zq50AjMkrWeLjjOR29HimwFpr7r3fIpVdYnA1fXctkE0oCjzdj28m/vIlg3U3GAIFyxQm1aaiSotPtyGA69DgYEi4D4IoBvoHUfzoX1N5KN7FCB2BflEZsFfn4TUEp
KbAWmvuvd8ilV1icDV9dy2QTSgKPN2Pbyb+8iWDdTcanNlkxUdZsEC86bV/CgKMzOBgSLgPgigG+gdR/OhfU3qr+LaXessR+mBo1j0OaoZEpsBaa+693yKVXWJwNX13L
ZBNKAo83Y9vJv7yJYN1NxusaCLyPrmo2tWiZRNBUTck4GBIuA+CKAb6B1H86F9TeFzdOw0akJzjPVpKANaPUOimwFpr7r3fIpVdYnA1fXctkE0oCjzdj28m/vIlg3U3G
ixuinOPSGN7ovKQEP1+RMjgYEi4D4IoBvoHUfzoX1N48kKWQPv4e9RRHkRiPX8hZKbAWmvuvd8ilV1icDV9dy2QTSgKPN2Pbyb+8iWDdTcaB3qTeKro2JOi503jolu6J
OBgSLgPgigG+gdR/OhfU3rqfar7vpoMpqEGf0T7aUzwpsBaa+693yKVXWJwNX13LZBNKAo83Y9vJv7yJYN1NxgpsB2z9oYJCSEUnhhi/rmU4GBIuA+CKAb6B1H86F9Te
M5G9xcGBPSyxmih0IG3lDymwFpr7r3fIpVdYnA1fXct7DdX1WnT/ZAUpg994pqS5w8xRG7h3qpFw/pnR02/rW/hi9MyMtWgVtHLHfL6R6jLKiCbRJr2HgYyrX3ljAm2I
KbAWmvuvd8ilV1icDV9dy2pkdgbISDlIhS1cURhpfy1EC1rAoVucQtTdo/IgWesZWQELFv5n8f2TNuPC2olLyEEAVVtqa6rqux1phTnwgeWJr1+Y0WAaMj/ktP30L3Ua
DMFHSJ0g+Da6RDne/AroYmrpFuo6r1bnqYAZKK/Vvyw0JT5HkplKokMNDrfdlZYG6s57HzcJ/ZMLsTIP3Mjj4CmwFpr7r3fIpVdYnA1fXcsMwUdInSD4NrpEOd78Cuhi
287pnpGpoG1LBDun9unJITQlPkeSmUqiQw0Ot92VlgbmfcwBd5EAEK07khe33AL7KbAWmvuvd8ilV1icDV9dywzBR0idIPg2ukQ53vwK6GL35dQLF8aNQiUMLhLLT3jG
NCU+R5KZSqJDDQ633ZWWBn+ogM0iQ0cv4IfXpLfA+xwpsBaa+693yKVXWJwNX13LDMFHSJ0g+Da6RDne/AroYj93vurf/0QfPWOCvQtgeDw0JT5HkplKokMNDrfdlZYG
SAMQj/WeMvD7L9v27IfNpimwFpr7r3fIpVdYnA1fXcsMwUdInSD4NrpEOd78Cuhi+Ns9g8S+AGnSGVoJ34gPJDQlPkeSmUqiQw0Ot92VlgbHtmrnQCMyStZ4uOM5Hb0e
KbAWmvuvd8ilV1icDV9dywzBR0idIPg2ukQ53vwK6GIAgXLFCbVpqJKi0+3IYDr0NCU+R5KZSqJDDQ633ZWWBko3sUIHYF+URmwV+fhNQSkpsBaa+693yKVXWJwNX13L
DMFHSJ0g+Da6RDne/AroYqc2WTFR1mwQLzptX8KAozM0JT5HkplKokMNDrfdlZYGqv4tpd6yxH6YGjWPQ5qhkSmwFpr7r3fIpVdYnA1fXcsMwUdInSD4NrpEOd78Cuhi
6xoIvI+uaja1aJlE0FRNyTQlPkeSmUqiQw0Ot92VlgYXN07DRqQnOM9WkoA1o9Q6KbAWmvuvd8ilV1icDV9dywzBR0idIPg2ukQ53vwK6GKLG6Kc49IY3ui8pAQ/X5Ey
NCU+R5KZSqJDDQ633ZWWBjyQpZA+/h71FEeRGI9fyFkpsBaa+693yKVXWJwNX13LDMFHSJ0g+Da6RDne/AroYoHepN4qujYk6LnTeOiW7ok0JT5HkplKokMNDrfdlZYG
up9qvu+mgymoQZ/RPtpTPCmwFpr7r3fIpVdYnA1fXcsMwUdInSD4NrpEOd78CuhiCmwHbP2hgkJIRSeGGL+uZTQlPkeSmUqiQw0Ot92VlgYzkb3FwYE9LLGaKHQgbeUP
KbAWmvuvd8ilV1icDV9dyzwC2FcfXQAeRWI3y+IIESZrHFUUG7jUqde3iFySOQtPWQELFv5n8f2TNuPC2olLyBK0Ycku/m6GH5G9648yFISJr1+Y0WAaMj/ktP30L3Ua
tG8akfbqhOO+2uDWwnIlvmscVRQbuNSp17eIXJI5C09ZAQsW/mfx/ZM248LaiUvIKKjV6T2lxsKTLKJs+DXpADqNafDcqTcpH1nyMYXOYoJz4WgPtkrwozxOaj2vEGe8
axxVFBu41KnXt4hckjkLT1kBCxb+Z/H9kzbjwtqJS8iNNrZKvgqMHVRvwzbsLwyzia9fmNFgGjI/5LT99C91Glhr8A4WbLv72AGL+QVM/m1rHFUUG7jUqde3iFySOQtP
WQELFv5n8f2TNuPC2olLyBgBr8b7x9sT3MiIU79WcfWJr1+Y0WAaMj/ktP30L3UauqYrqERkNHKnxP8+dhgh7mscVRQbuNSp17eIXJI5C09ZAQsW/mfx/ZM248LaiUvI
5QudvoRbr9yVEifrkBs8zYmvX5jRYBoyP+S0/fQvdRqb0IiBU3dP/d2SgCMxE3XoaxxVFBu41KnXt4hckjkLT1kBCxb+Z/H9kzbjwtqJS8j3hvH8w1iIpPVJPMPOP0Jv
ia9fmNFgGjI/5LT99C91GjTT7PLL65fLvB0aQXjigx1rHFUUG7jUqde3iFySOQtPWQELFv5n8f2TNuPC2olLyPfcQr2OdOkGi0NueUV6w9aJr1+Y0WAaMj/ktP30L3Ua
7dFLIKxLZ9aFK435RQ3k/WscVRQbuNSp17eIXJI5C09ZAQsW/mfx/ZM248LaiUvIsTYH8hjduyw84J3+KiobqYmvX5jRYBoyP+S0/fQvdRrpgAUBscjqnUk+2mqpl3Q2
axxVFBu41KnXt4hckjkLT1kBCxb+Z/H9kzbjwtqJS8g2HwmHqzVPY7XRyjNT4pJUia9fmNFgGjI/5LT99C91GlP1LbcEKnYgw3SVKHJw4m5rHFUUG7jUqde3iFySOQtP
WQELFv5n8f2TNuPC2olLyDxYkh7zMd/QgNfU2oJ3RYeJr1+Y0WAaMj/ktP30L3Ua8zRr7+81Im0rS7YFZP8mrGscVRQbuNSp17eIXJI5C09ZAQsW/mfx/ZM248LaiUvI
zE3AKDkKMayBxXb+Ld33aImvX5jRYBoyP+S0/fQvdRr6qwOFGgrUkGh3lG5l7u8JaxxVFBu41KnXt4hckjkLT1kBCxb+Z/H9kzbjwtqJS8hmNHDi1kALfVvr6f/KZJic
ia9fmNFgGjI/5LT99C91Gout9b9U4bzqhbpwFbTQ/GtrHFUUG7jUqde3iFySOQtPWQELFv5n8f2TNuPC2olLyBNx+jk5grmg+qAeOPvzmemJr1+Y0WAaMj/ktP30L3Ua
hTseZjaETGV2/gqEOTVEVGscVRQbuNSp17eIXJI5C08bdr5Rw4nwbjrFH2dX+O7NbhT0JmX44iFIMrJJvh1k5ImvX5jRYBoyP+S0/fQvdRqrB62rmN5xStal3qmZ5QZW
axxVFBu41KnXt4hckjkLTxt2vlHDifBuOsUfZ1f47s12CWSZOfnxWxsv7PUUFftmia9fmNFgGjI/5LT99C91GotEgQ8e07tm88ELew8CHs5bGhXGINzfUvGWs/DYIhlf
h0PTKiurs4pFAGcS7dEimcqIJtEmvYeBjKtfeWMCbYgpsBaa+693yKVXWJwNX13LsBXjSSPfNUy436EjruMyeCqPZvSsJfn1fRBz/Evb+4r6gj/hPWpzJSMgZ2rvq5p1
yogm0Sa9h4GMq195YwJtiH18CNVEugvM7D4IfFS+oqtpKajDTmtl30AI8XzTfgSYF3aQQcZrXtDdNulRFhZ95Dg57Z6VZShpm+zbva8NQvr7rICpy6vrQuFpgCGDT3b1
rn6+6YWNcZ6mkpF4B9S7++7V6+pQ7z2ofAGj+ruE9xfKiCbRJr2HgYyrX3ljAm2Ig3EXTn58wwiGNPL7MS7te4jbIZ7ACAdFU2Qs77QgQLhyO94DM77/tTnxjBLslRoX
XdlpFSC9+YVc0iaFRxSG//foKSoEtXAbz0dSQqNz7gAykjPpSkhcwQj/OydYo4rV0yGRnPZE1s62DA8g752IHP0NwjVoPQpcuqk5KJIg11hyKFIWQEE6a58j+AkMv7ic
i2WtS347aixe0KbQSsWojcmYlOeADlxWcAPrGWSW0F6WYnCpLHNzGAC4XS62ftEe3gRHoQ0bubQUMPVuAEVMOtwPx0FAGBxmMHPXripzH/yzcoepBOgwzgCawSN/z+bR
KbYhdNiWjh8peKQdr+s8ajMQfksFkJQxB3BebIhcd9cf2JiOmqgDz77PlYWnpGaRyogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YW/d4ucwAkikPsRv6s1HcdV
OAWTZCKXz7wIbENXZJosNVIA/02+6sVA9jyIA/xPGUox60vdzazTWl9AlpLjoud6yogm0Sa9h4GMq195YwJtiHRDKVZNP4lSwf13PICjvgMkCVI3QfLkZlhMZvFqxXcB
fqU0ivsk3q9nShpikBsQ2aqvRlMQEgk0zpj9ytY4TNFBVGvT9cNxscOK2hBOJXKUyogm0Sa9h4GMq195YwJtiPa7MB+UZd1JHic/n+t60++uLUiaGSbRvMiO2Y5sCASN
zTueu9UaKrMaHCXH6TsqHKk+HwqbFIiNduUhYkgNDzbSQXL2m9w9gHqvDLTrcjziyogm0Sa9h4GMq195YwJtiIEayJwYGQ9fRzfY+QWc56NWipiTLetluFwCQyV1q4yS
DH2RdZ2YNaP7I7sYFZEz4Q6Om/thnDZey2EFlRJHzBLUAJinUOekvV0p2S99ct3myogm0Sa9h4GMq195YwJtiJ5DxCzEkASNymFUZ4DxMUYTiY/nIHLUaG7nhQ7jQlgh
s4d9zeeKhfMMXKFEPYZc065+vumFjXGeppKReAfUu/v3WxEf761t7i+hMnhJ7Sg9yogm0Sa9h4GMq195YwJtiINxF05+fMMIhjTy+zEu7XtUgg6xaVOo6C2dhYizYT38
ikcc94OyHr5c7PXMMHznRl3ZaRUgvfmFXNImhUcUhv/92zJDvpW1dUkdbWMunoR8Ms6Yp83sbEijSPVFltsRMNMhkZz2RNbOtgwPIO+diBzzSzW7Y6odhObQV3/Yyn/o
3ea9yDxSSJF3wt1QQcMeY4tlrUt+O2osXtCm0ErFqI03nTkJetDTBC2uEW6f6gB1Ms6Yp83sbEijSPVFltsRMN4ER6ENG7m0FDD1bgBFTDrcD8dBQBgcZjBz164qcx/8
rKjhvONqFIGWIfPho+7gcCm2IXTYlo4fKXikHa/rPGpRAR54d8OD+g/ftfkcL8wqTE+opLm2tAq76/ZYyqpnPsqIJtEmvYeBjKtfeWMCbYhtzH0Dd64lp9Q9mHuXW9mF
5fboCS0G6zJmeRqBuyulPaBEq5qlBjM6tRS0ezL84dSoGd8+DQae7WrPOwePZ/KN3MH3yNHRPOMmuAV3JC21M8qIJtEmvYeBjKtfeWMCbYh0QylWTT+JUsH9dzyAo74D
3h64Z5Vt974GrBSTvC73oA9Rw/+S5UHfjJdWkfIeInSqr0ZTEBIJNM6Y/crWOEzRbztmR78bGJkkrUx+KGBxj933cmDSk9SKNleh+t8ICqFAyaqwkAgzq4ApJkwTRqQM
G56S0vu8OQOPhzMAs60hlkmV3UcDeLGhA/7PNcP63UygAO89LggsGPT91VUubNtR2IxgPx4X0/eBdEw8eySRiMqIJtEmvYeBjKtfeWMCbYiBGsicGBkPX0c32PkFnOej
AIgEYrDm72pdPGqSWEl8rzTOYSt5l6buY5IsJUVrGMcOjpv7YZw2XsthBZUSR8wSbU9Ub95AzUy2zeLfcaiG2pvTPN2jZrtsTg11onp4vGwssSL+kQiAxhrtE5GaNEr0
qJI7YEbeIAYkNBFAqjXCBKowGgD7cb63+1hbVEofIyaufr7phY1xnqaSkXgH1Lv76L+E7lZtFVHIJdIvKyg2CqZq0xwMNhJ3pNNT1vrO6bBx2TL+lY4mzdRBmqXHNKXG
JDqsLJwI+62VjXfg0kQlU0ZSqlQ17xDj9ZOb5xF9CRdd2WkVIL35hVzSJoVHFIb/9+gpKgS1cBvPR1JCo3PuAD/aqxE+nhezx+L6LFdldSeyfwRwZreucj+evpHCy9wX
kjcNPXBp4PFAtM7mq3J81RgVNrLtYur5z3hC6MV41fOLZa1LfjtqLF7QptBKxaiNPFXdVbtxFepJZP66g/nVKqKLpsBWu8O/ayZjdJtoSjXedGbxxIYjJ7I/1TyTy+3O
K09CAaC+GdPoTocIAxv5eF4wFMarttComGaQ3L95DcFuJ7T/5M0cUlAxtp1zhkMo4buRwVhLdfLrgVnZx9I2k0zWsPoOd0KUSX8SlgtD8MvQZueJC7GqmVyxhdkNqLPc
EkaolafW3+oauiKYwUAYVpzJPIvrIemSLOsF+r17NbrjWlyXc1Cu14KZoFwgI3/GSiGdAIboKY9SXPzUKSG4Wxto1TruR4eZ1tECV23cD27cWjM3yyRwaD6xLOY8qz3h
FdJkT329i7COnhM1KYxKoewAXfTS2aPIj4vaTjjhAnZL02u6/egN6rk+L/XAaWWNqq9GUxASCTTOmP3K1jhM0W87Zke/GxiZJK1MfihgcY8A4AEl4pNNCx46HLNELETD
QMmqsJAIM6uAKSZME0akDNScD1CgcTMtq9SDZI3h6qM1uJcjBHPTnQWALUhXdH30qT4fCpsUiI125SFiSA0PNq3F75sspHOCwJ64J6v6T1KEBLLZ1EW6iGDgQldTtneC
EAR/jjP8ddXOJ3kaq7u1rgCIBGKw5u9qXTxqklhJfK9VgaqGdoEGWCj2DJ8Cyi48Do6b+2GcNl7LYQWVEkfMEm1PVG/eQM1Mts3i33Gohto3APUooeWprIyvWDqn4w0X
9aLTJYYjqbMSmwTo9BxRxqiSO2BG3iAGJDQRQKo1wgQTI5xsXBexaA+GrI8a89h6rn6+6YWNcZ6mkpF4B9S7++i/hO5WbRVRyCXSLysoNgogxH19CX5f9PM2RtDSwyUv
kayhKx59LtadPcYnbadTwiQ6rCycCPutlY134NJEJVNiTTMfKElmKfajDXBc1z+1XdlpFSC9+YVc0iaFRxSG//foKSoEtXAbz0dSQqNz7gA/2qsRPp4Xs8fi+ixXZXUn
IocEr3+XBfL+Ds8ts3lrTpI3DT1waeDxQLTO5qtyfNVYCRXYlweMYlnAMqeOqmB/i2WtS347aixe0KbQSsWojTxV3VW7cRXqSWT+uoP51SrzPzlfeAXuh7hlNmd9G8t2
3gRHoQ0bubQUMPVuAEVMOitPQgGgvhnT6E6HCAMb+XjHngGjHEmQVrUpEhq/RPI6+ykV3+CGzMCsZ5mBvXObHsqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiG3MfQN3riWn1D2Ye5db2YVzOiHGZV6fLwKbnZqpEGRo8kItuzEWqMjeJeBS026F2kohnQCG6CmPUlz81CkhuFvHfWojvrM/wXvjC8LipbjA
NtvxKKotmzizr6EdreqNIBXSZE99vYuwjp4TNSmMSqENg2ydJdNhjlLcGNXUFOTlromS5z4xoabrn/f140I9QqqvRlMQEgk0zpj9ytY4TNErHOuN78XnBTUn0bW9m91f
3OI5gbPyhZM8tN9nD6LOHEDJqrCQCDOrgCkmTBNGpAzVUnlsNHW4rXRwkYy/wmKjQSztJjqLeQ5+k/JCMA/RBqk+HwqbFIiNduUhYkgNDzatxe+bLKRzgsCeuCer+k9S
17QSLqNva2UCN9B0/Z7NJXfEe8VdIKb3hCk1MFzH2153aByBiKdJV7+dZ6QR0Q05UUJQv7vYyr/E6SFviQIXyA6Om/thnDZey2EFlRJHzBJtT1Rv3kDNTLbN4t9xqIba
BqYPlpGmZU6AkbsKQ6IOdbyFAbOwJZE3VTubHW2Ne3Y2O70I/6fuuGkGRLal6DGOf5aHbAbHKqnTwG0JFxkMqK5+vumFjXGeppKReAfUu/vov4TuVm0VUcgl0i8rKDYK
I6r9hTz9xeBBxqCPNQs1FZ+U9AFUZdQiWBYPycKk3HEKmF4NFJvGK2AMp4SLhywInBNeLnLBAvtZQr53wNoDkV3ZaRUgvfmFXNImhUcUhv/36CkqBLVwG89HUkKjc+4A
RNvQ9yRxrJMSFA9jFrgR8FV1+o51qocFDgp4YmKiDuOSNw09cGng8UC0zuarcnzV7mfcNI2NA6Tjd2u7J8lL04tlrUt+O2osXtCm0ErFqI08Vd1Vu3EV6klk/rqD+dUq
ooelsXGfLkOi9pPYGauRLJKRUFZmYkQzT2BpWwPU1bcrT0IBoL4Z0+hOhwgDG/l4+layRTwpQrR1P7aBFUbLCmGWIGb9SBiUgm2ZK1PcxgPhu5HBWEt18uuBWdnH0jaT
ehxJh26eG0iu/A7AE000wK4FvBR3FaZW5+dshhRZ4MISRqiVp9bf6hq6IpjBQBhWESK6pPhS0GtLhRevlu/V7ByANaqg5+XEI8TTnyyIqmZKIZ0Ahugpj1Jc/NQpIbhb
x31qI76zP8F74wvC4qW4wGCsLHAk1MQktW4qfSx95msV0mRPfb2LsI6eEzUpjEqhDYNsnSXTYY5S3BjV1BTk5U7O46rzohS2Te9owVgqkeOqr0ZTEBIJNM6Y/crWOEzR
Kxzrje/F5wU1J9G1vZvdX+o5Ku7pdapgY3tptCa4V5ulJshuvalJyhHArIhh5o9U1VJ5bDR1uK10cJGMv8Jio6eZwaTSYiJtt8bLya9VOwCpPh8KmxSIjXblIWJIDQ82
rcXvmyykc4LAnrgnq/pPUi1vTiswGXIcxTi5U5jWEvx9SChKNknSZ8s69N+tqhXOxAAo/hDCFF4NQ+yjGK31QcqIJtEmvYeBjKtfeWMCbYipUeA0g95VzZWmFRXXU//A
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYieQ8QsxJAEjcphVGeA8TFGGFPZhjO0p9AR9Gt4g4m38ic/zDhU8lPwC5MfkEe7Zzp7BEIhGZ31+yYfbzxoBQY6
LmKRiI2lIu7X97POMWrj68qIJtEmvYeBjKtfeWMCbYh+yGZrmBneblZRmw9FMfTXB63wui7SL8kGXa57GDgbl5JOvdX02oAhGWjxZAYVa7m+Nm9RcNlplZxzYEIyhLbv
CnErUe9Talc1aFyPDA2mlMswjVqqyFe8TfBKizBIh7sPUcP/kuVB34yXVpHyHiJ0qq9GUxASCTTOmP3K1jhM0Ssc643vxecFNSfRtb2b3V8r25FgHUwak/Y52YK/nCVY
88JKhJEpeOwRxLuj4ic/RfXgIbG2KXL7lT6fOiJjyKrNIuz5P/6n+zU0W4Q3q6kxsVKQRByGDQIIrBrQWW+c6g6Om/thnDZey2EFlRJHzBJtT1Rv3kDNTLbN4t9xqIba
HFPlYW04EDnCYxWJ7hWMx1wXhBj9h8A7jdM2yQpq9Sb2hNJkUWtvcXHVF4k+rERCUAwbLiqqh0viIfFExnoOCgeHAGKR1sKCOTUp54XcaBBd2WkVIL35hVzSJoVHFIb/
9+gpKgS1cBvPR1JCo3PuAI6jjeD/oybZXurF3QEUExPtiu0zeJm4i3gWWCB8RyRUTX90VAj5s2hN0DcK1cpi9HfhVAV2dy9zisaodInfmAyhoQQYmzpGWA5C+VnN3r0U
KbYhdNiWjh8peKQdr+s8auG7kcFYS3Xy64FZ2cfSNpOiDFeTGUmz2p2f9KodTz4YtkfY1LJl/1ulAgVsqliNiY3l1ow3ID6NyfDYYSmbMV2Jr1+Y0WAaMj/ktP30L3Ua
redv9QPpHaMI/dmeM9i511LTkzuz3QSGh+F5Ij2Hzxr4sYtYSRTxWZaOX6vJ05Yjyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
9eAhsbYpcvuVPp86ImPIqlisWByskj5/vDXqZLmdpn/utGKWGv+cQhDubKk0VgnODo6b+2GcNl7LYQWVEkfMEm1PVG/eQM1Mts3i33GohtocU+VhbTgQOcJjFYnuFYzH
75hDSmaNh1GI59Ls6CRU4NkXW0QWBVb6JsOzT7pVheSa0pY/DuluUIHvmvQa47tUOP8FoDq0i1xV19PKzLcyqd00NeWoIXHVF9/FAs6jOM7KiCbRJr2HgYyrX3ljAm2I
yogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2Id+FUBXZ3L3OKxqh0id+YDKbHhnupiXh7Cwqipg1XPfAptiF02JaOHyl4pB2v6zxq
4buRwVhLdfLrgVnZx9I2k6IMV5MZSbPanZ/0qh1PPhi2R9jUsmX/W6UCBWyqWI2JVcSGb1e7nDfmH+SghWf0Cf9aBBcd208zZRgilk09ksCLRIEPHtO7ZvPBC3sPAh7O
Jo30qpEowBX7YeLA48u0/Vi7RZftaIQzxdKJ+LTfsT/KiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYj14CGxtily+5U+nzoiY8iq
8xb0gN1Y/6WnfBIMWnFjF75GC1/5ojCuIkaaOCknpFfylwJgiF4ltfD4OAp4D1reyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2I
0bs3uyhPJXfV4SVgiJm4yA4u8YGQBgcJMkkXD57lfIOYaRMyMkJ8oCQ+qFOTVPDl6tDCLQ++zkMZWMRtcsNkQcW+v893AwXKS2So7mgMfcf7ZigYx3D/J/uOoduvkkLO
imwCyuUgSJzdNdWn1mcBysN4xfXnrZS8v/num2K0qNjefW2JWm2UOly4NhY2h/B9EmbJi1qURa6f1x8gsCQYvl/EPZBLsSaFqRyddkA7EIe9ZNFLaV9ubOG0KtM5rHpq
nNS9RrFvHHpV/gNbiDMtXBWhaW/3HwJwNJ5QOXIwwPL0T/g7chVMi+ILuIUWEUQPwkjoIJewTh9jGdn99+Kgw7l9zi1VkrD9kTvfOPLI4QbKlNzlprxvnTHOpMJ7phpz
5zbe2d1YIJhmBuZnAg6erFdLvf3DL/HvUruzy1Z3NWkRlBoHs+ToItjtsiNX3p4usMFN4PESh/NljSRIa0+tFFI2M/a4ix/D3PRGRUGP5susYSXhlSEO1LgUYU2nhj6C
bDnXjMPiOdR65htcTFryqPKdhQTe0sz1UxiGLzU/u2Zb0A+O/j2+WWIKyZo9yoMjcAuWgUz+zCHqd7/yuQAS2tt8hy2pwr37UeY8AMqLxYcAGq2JHUVW9QOebExOUww3
VB9PeGb+j+CrtZnzFEW/USStj6YIp9+YhlSQo1sl4AJJLB7KTTf2Uj3NGrJWG0azxt7ussSBZ+P/RYoOY8YgihK1zpsX3RaKxD0CyHxUjn1MCHBT9YSlLpfO4Prm8Dmk
rPGsGD4oSGGu8vrZ2e4bejX6nd6mKDhUrO1E/iuetdkbsrSFnOqFWlr3z+m69YNRQw+8jHVTe+rKoA+dMh5IUTWAupfxYFLfGXNEynfAQPYnUtKcVL0y166x5QYzBQwr
cdeRDbFoGyCsHFT0nIKUj88Jk+00ba7AyGakdPek1NeMI9VW6hHSIsjzcHkL1Tlnm7OUpyqr9qjffPe27Ox6Ap8aY2klu4tCPTqozyajDuPAq1MfG7ua4ommDuLe2+U4
xNLkLvGTfBmDplhgusYrdLniZSs2iCi7ZeesRoIQJFSbs5SnKqv2qN9897bs7HoCnxpjaSW7i0I9OqjPJqMO46djWfJViXW9BU9Vx4jdeQjE0uQu8ZN8GYOmWGC6xit0
fvlpS+vpSmNu4ld+HTVI712wnlmOiVIwYggkI4iCRgjeBH+xjaMs/mxQh2WrrCdr068EDie5dc1eZx7ync01BQ/ip26VSFsAuui+BFHynu3N2zbtICS7LPpyY3GIS8JX
X7ZnrmaR8F21yRQl7ZH1B01Lyl97mJGwt6YosKrRCWiD7tbtlAz0oyO0X1hnxpHL8RO4MPymqrwFvU81rUqGFM3bNu0gJLss+nJjcYhLwldftmeuZpHwXbXJFCXtkfUH
5XAuFgG4iEmOklgQqTryk4KxX1sXKQe87JroI3esbqVbrMW/ubdG5dqi54/LPTjujWaZstcOJ1Fy973DzJXAZ/RP+DtyFUyL4gu4hRYRRA/YO869ra5635LE2wAhdoI6
zBaBQxdZNXNj3vNOVzrQrTXq68RJ+GR3kh63pfTu/eu7xxsPXIb+C3bTmbbqysguGLZ5c/vV0nbjrM5QtVzIV3uwJIUG7kQFXcV3BLttfx+X2qTQdbIyrf/YJe6eN0Rk
c5URdJc9QHbnn7lifqez3YXE+8h2lsqIY/KBOl3iAOdz2qej5sV1BXImIa+YIhe36jc3ZSNOaJVzCME/QMqZ4hi2eXP71dJ246zOULVcyFfZYxH+Aaha3CSV26e8ak7C
UjYz9riLH8Pc9EZFQY/my9DesKTryjSyqDAvUC4nufg0Aua0RvAFE7Sf+NwlnYvdOWAFTO79GREGnUVL/1bKc4sHOUlVxDcR2vy+5qhE9yxtctBl8xEzZ9ui0Y24f085
aD1nqpobrx6GDwS9FBMwXVNOWd0IUBqrgzvKmtZDJ43MDqkq4eKg2UajPIxLsizNGLZ5c/vV0nbjrM5QtVzIVxacA9EuDwC0IM/cvTM2WrH0T/g7chVMi+ILuIUWEUQP
vV+pOgiIxWYywnpsZCm8JJ1xwJEK7CiHmuBKgnWzmUcs+w/c5ew7L1IeI0mFvBrbEcROy7CcihmDbhrXtn6xLH43+xsJ20+8V9fnCRh+9l5oPWeqmhuvHoYPBL0UEzBd
+mishkReL3f6IUn38AACtnodGXGW63vD2Py1zBG77AnCWDBqG3U/rAyKc4PZdDKQ3ucRhIS84X5SJSfa1o87xvRP+DtyFUyL4gu4hRYRRA8uoQpj1uSHnxbmcMW9F0XW
hcT7yHaWyohj8oE6XeIA56U0Fr3oLJPpwXs+eklXZnyve4VXL4QomSBdP7zg6hRwCHDfHnr25ZcUlOdQI6wlBVmKBtkMoN013XNxh7tjOhYCtEWOlbO8y8N9vPzmIpWl
8Qim2XE22j45hy2JZADfWRi2eXP71dJ246zOULVcyFf2GlMeUjzXsw+kaPoRQJfVWlZoQFVdXWRDqQKGCHhB/zaq3BgHmRMWDzkRvpWiqEkFZLbYbt7YCrbWWdqEXKEB
Kl4HuRgOMcuvfYBonmmyPT0Y2h3Rt5WJF/BpT8mVQcxRiR9Fhkv0ZwVKldnKpzCYj2CwAxDJyf1zGs9O8LPH52BvlKgyjuOJ6qb0TJeiJQ3CWDBqG3U/rAyKc4PZdDKQ
f3t0z45lXYabZniV07P2d1LvzXILZF6ZBj4xpTeZd7RvJrk4BotvYSssLfG82ljSUYkfRYZL9GcFSpXZyqcwmACaXVrnZ96gS8W8iYiKLX0sDU5oLp2YZwkEzEDl6/pF
eLHBzQPhOSax+GnQxQVR/XTWpN5BrXuNJZpEVhJKG9CkO1Pbzl4V8W93GuxefVkFBH/8bwTsbWDiBRks2IWn/3N/Bm37uZHniDH0S6MFMrUw0469cnrjOubhMN5rTW69
fl1l9+qa+UiCIgnuji9c+HnzUtHX/nMF3JGSzByeeolRiR9Fhkv0ZwVKldnKpzCYN8jt8G5dmVl5z2VkBEHmBPZJPHVeUf/C/PSIkzr+cOgIcN8eevbllxSU51AjrCUF
X4RQscDfrERbv7VGPOSaZ7sOkpB1n/9E4jfOlTDFDLjbifQkoF64pp1DcET+cy6Hc38Gbfu5keeIMfRLowUytZWwd6L9NXzOQhn845+Kku/OxDvP4PbsLKiDIawSBsIu
Sn4B9/eVbnFc+7d2ZruzyaygdwYa4nzjiQnp/QNflSapMsAFZpquGKx9lKye6R7l+3OHWJSaHNrxHdOFC6DtXMJYMGobdT+sDIpzg9l0MpAvU4Ckgfo3b2I34Rr7sRMc
hktDTRqnq7W6Cg+SeAjI1xx76XmdxllsAL23+ls7OTu8LvUypHyymatYyzHl9SX8RalIwPKNbhDswuP6723RpOywbwQnC8lbVu5G8VqCgHL+JWiTUS2mV5zTUL2v0xZq
DUVInKTnm4eoMZ6evsdxBgG2T+EcNWw8LDpebz5p8itL1YmSsXqk8Eo46l+keG453CESd8FHfUYRJzBwZYcOE6GYk8lgjnYDP4RrARAe+g2ZLM7CPlC8j2jO2rLwVsbp
sXpnoVzyEUzAZ+bg9Unagrl+sRZr7sdNyMquWoIyKpOpPh8KmxSIjXblIWJIDQ82rcXvmyykc4LAnrgnq/pPUj64+JVA8SAPwyc05tHZm3FT2WR+q35TTk23PdmsQjA8
O3k4rcxAoNsVtXkz68BTisW+v893AwXKS2So7mgMfcfxH6Y/dnI3TKHHWFadlBxK+Gz1HcG3zSZn7HE59S8LgEIMEOKNSg1JInKKzeN3rhZZAQsW/mfx/ZM248LaiUvI
vseOISzfypxPQeNwf8vVk7BLB29zX0yznPwExGGjxGojPlTJc+aE7PSzruqztFxmkq387EtQAfhUaj3utHaDDuG7kcFYS3Xy64FZ2cfSNpNM1rD6DndClEl/EpYLQ/DL
oE5XJsc5xWskbWNhzI1R3YXS8tvV7KBA+CbFCuG96No7eTitzECg2xW1eTPrwFOKxb6/z3cDBcpLZKjuaAx9x14wFMarttComGaQ3L95DcERt3F9MrLiZrH5ZSsud7qL
PeoiJVFrjLUV1sBGHWbzOaqvRlMQEgk0zpj9ytY4TNFvO2ZHvxsYmSStTH4oYHGPXwm9cRqMAUECucGniPrFKDtpGIfLICEFMPRsoxGgUnb+uqpTYb598Cau/itPQYiP
xrqlDRFDM4VekkAFoPghdYKWQUszSgTV3K2lhiUTnSdPn0SV3FwP69HfRqPl7u4uFgPpaMN0R/oDv9yk4m5Diq0hUEoRF27QUbMYqJZ+6LXov4TuVm0VUcgl0i8rKDYK
5lrzQRK/vccZo2cGPda8ZMPMtpWKcnwbyq26sOhxeriBP0dUDkM1hct6UAILUDvGqq9GUxASCTTOmP3K1jhM0W87Zke/GxiZJK1MfihgcY/MJz0rlvsouiABJOuHTCN2
dml+IKrdOrbVOL2fPuyext0teUbdk1LIaoMoUFgIPMaze6G5LTlpIP6cwQ9HIOPV7ABd9NLZo8iPi9pOOOECdsTz89aY59ArpfwCw3gWA1HuQT9rPM44y+3yD0INerKj
AbZP4Rw1bDwsOl5vPmnyK21PVG/eQM1Mts3i33GohtrM3po67117uHQTB8F+Bdb4eBqpBnXMz/dIW2ybx7LJb7wWL+C+JlSTpdhsSNRe8NZwIPdgr0N25FAyGdBWDIlJ
NA2wTCemsw/ciANN3xf19JllE6m+ByMl91vJza/j3LepPh8KmxSIjXblIWJIDQ82rcXvmyykc4LAnrgnq/pPUtF+wTLo59r7D//4LTly2ovEXHUf2z4IMrQYommpoUfq
xrqlDRFDM4VekkAFoPghdYKWQUszSgTV3K2lhiUTnSdrJUcEpEPj53yuROW1yILSqT4fCpsUiI125SFiSA0PNq3F75sspHOCwJ64J6v6T1JfAOXTng+tyQchEWSvfkh+
CZvM8TFuFCkCBNGL9KqPICibGYWYAWLJ046Rr/CXzi2ze6G5LTlpIP6cwQ9HIOPVxYZICqBGtB6VVnOsjp6s7jRNCkq3gntxNd+H3bJfU5Y8Vd1Vu3EV6klk/rqD+dUq
Y0JYOiEKnJ87yKwKyhG8fPVuOwDEFXd6lqvrNNFmpi5VQ+4YD+qikOjYLhDAPd63H3ipDgvurEl+pLsnNqENB8TCiPKQ07B0wAGGvUcu2pvdlhcbDJw1qzPe+6lBg/4t
2EpW37RyZj6ORbsFec3PxwmbzPExbhQpAgTRi/SqjyBtTPWnx7UUPmw0NSR1DvXlWQELFv5n8f2TNuPC2olLyISxRLLkotOaSGc8as7ZX/H+VkEl4sUJJyTroob1/JRR
DM4Vsrz2Dm13VDwPxjLfjikjxD7yEsRy6in036EogDT6TKnsRDdUgZETqEJiDdrMSpeE2x6uLvShqm2Qy35+40ohnQCG6CmPUlz81CkhuFtdkVJCCDZiGdxvGp4yaesw
GDMHPlgIp+vVE9oh6c9WyQ8K4ZpMDUn87sv6YKij6Ejov4TuVm0VUcgl0i8rKDYKa7GqFblDC8hKFcSB448kIFymXaZV1Swl1y1luj5g1NExIaNyNYfe8ZzGvK/qK3/D
McSWsKWAChUzquZEtP3a10wJBwth9hirsiG83G0F4ECCepKn2NgEZy7mYul1Oe5g+PB8w2FAcSpQL6H5xGQkTAfpMlyT2iYxIV1YHSC5XAqAvn1wjCzg4scitxorJ5pJ
9+gpKgS1cBvPR1JCo3PuANXaCyx9L6aNc6X04tVIW00FclMUWSiAFf6ix+h5ZP+NqT4fCpsUiI125SFiSA0PNq3F75sspHOCwJ64J6v6T1LXtBIuo29rZQI30HT9ns0l
cH5hYGsrLR0gIfubVGUWO8a6pQ0RQzOFXpJABaD4IXX2X6tOzAKTwny8W4ZPyUuHbYdKmI/2nCj/XGGOTKzgoqk+HwqbFIiNduUhYkgNDzatxe+bLKRzgsCeuCer+k9S
jXyBcO7TeIELGCUj1T1K0IC+fXCMLODixyK3Gisnmkn36CkqBLVwG89HUkKjc+4A1doLLH0vpo1zpfTi1UhbTUK8TSSTPP+sNxpmIcPGHx+qr0ZTEBIJNM6Y/crWOEzR
Kxzrje/F5wU1J9G1vZvdX/UzScAn/MLBl4JLApLGWIEG28dc5pM2iGe3Ybje4nk9fv3Gij/pC7X3nzbuBUF/7/ce+Eulog6JJlIGxSraKS8I8FHIYjTdNWg1SIti+L75
qq9GUxASCTTOmP3K1jhM0Ssc643vxecFNSfRtb2b3V9fCb1xGowBQQK5waeI+sUogL59cIws4OLHIrcaKyeaSffoKSoEtXAbz0dSQqNz7gDV2gssfS+mjXOl9OLVSFtN
c52Q6sLbt/UaGxd+a0KrD6qvRlMQEgk0zpj9ytY4TNErHOuN78XnBTUn0bW9m91fDx7EmTZqu/JlLjaPUFAuXgbbx1zmkzaIZ7dhuN7ieT1+/caKP+kLtfefNu4FQX/v
9x74S6WiDokmUgbFKtopLykzZe7vxfgXqEkZvZfHkBqqr0ZTEBIJNM6Y/crWOEzRKxzrje/F5wU1J9G1vZvdX8z9jnGrm0CzGA8gTq1iTtmAvn1wjCzg4scitxorJ5pJ
9+gpKgS1cBvPR1JCo3PuANXaCyx9L6aNc6X04tVIW00SQaRIyKxrkdCK7Hb3jOfSH3ipDgvurEl+pLsnNqENB99VD94fkvjyTq5So3V+89tJ8GXh26rvWrSK1X1CqgXu
/8e5O6dA/S1VpEGIiz7CLcW+v893AwXKS2So7mgMfccSLB/l458jxkoBRJu/27NvbhiL0b4PpSmBWKYtOKEtTjEho3I1h97xnMa8r+orf8MlQS2PNBF3vBJ9uhYc/8HY
+nL6D8FishjbN4eqaykLxh/xQiG/RSzPesEBU4357KltT1Rv3kDNTLbN4t9xqIba6meb7u1Zm39a6kjbNv9Z8yT3ec3Op6uZ2a2ime3z7DsxIaNyNYfe8ZzGvK/qK3/D
JUEtjzQRd7wSfboWHP/B2LDZDHhIHcaZP/RoXPkQVef2Lh3Q0PqsdHaISRidckeq3WiaDqn4WksMQqAppsVSuR94qQ4L7qxJfqS7JzahDQfEwojykNOwdMABhr1HLtqb
hC+yCArTdzetdSrER31G79XFT/CjC/3fZmqWejloixrGuqUNEUMzhV6SQAWg+CF19l+rTswCk8J8vFuGT8lLh0wpgwgDy3TyB4H9zIv2D4qpPh8KmxSIjXblIWJIDQ82
rcXvmyykc4LAnrgnq/pPUpCKw65fAh2KZZAh9z+qqfaCepKn2NgEZy7mYul1Oe5g+PB8w2FAcSpQL6H5xGQkTImmK9pDAjMymiSgvIZbnu2Wlf2N6lXDvwVmgCsPGLCT
/8e5O6dA/S1VpEGIiz7CLcW+v893AwXKS2So7mgMfcf7ZigYx3D/J/uOoduvkkLO57FTCVkhR74Isuq3UP3BodebgFspf4T/qNhOPIaW1NZZAQsW/mfx/ZM248LaiUvI
hLFEsuSi05pIZzxqztlf8dL0NyUqqmPT+HEKPWivr2leFNkyAoA0POwH52nmvWdiMSGjcjWH3vGcxryv6it/wzHElrClgAoVM6rmRLT92tf5H18vvwqVg3IKV5ivs3ik
qRxZ+w2BPjFCMWe4RxvF1v3ZpKz0cygtR6mhkfDEe+EYQbNd35207eMsb/CQucCyWQELFv5n8f2TNuPC2olLyISxRLLkotOaSGc8as7ZX/HS9DclKqpj0/hxCj1or69p
W5XAmUoey8ZR15z3OAnz44XdpGqHOoNlnsGGUGAp7mzURP77o7LEoIJWlhQcvm27xb6/z3cDBcpLZKjuaAx9x/tmKBjHcP8n+46h26+SQs6KbALK5SBInN011afWZwHK
4xUtcxn+6lqmD22gyfcUr8E5Xkxu8HutaJbbLpv25E8xIaNyNYfe8ZzGvK/qK3/DMcSWsKWAChUzquZEtP3a1/kfXy+/CpWDcgpXmK+zeKQf6xWa8wqk0AR+esHtnsIZ
OgUSFjMbpE1FGNOp3sN8E0ohnQCG6CmPUlz81CkhuFtdkVJCCDZiGdxvGp4yaeswEsQZI1smfWMLNvbttwQXB1+g+ahR9MomsztQdwoKfHsxikWQ0JFi0u9kRTfjtBLb
8Cvc0BOUKYs9tGWaK2Q9+ui/hO5WbRVRyCXSLysoNgqf1b4ms4jHm2DlgudsQFsNZ9mVT7SVRohCNCuzwokqwh1An/A3kX0V+/iGMAKq7ThZAQsW/mfx/ZM248LaiUvI
hLFEsuSi05pIZzxqztlf8dL0NyUqqmPT+HEKPWivr2lblcCZSh7LxlHXnPc4CfPjlApwKh3AUPbY8/7BfiK+VoC+fXCMLODixyK3Gisnmkn36CkqBLVwG89HUkKjc+4A
jqON4P+jJtle6sXdARQTE/tQfx02f8/IPBfmkDiknVCUXxDj1sgNV2SZvRrDpvPDBAJHag6xO3rs1E2PghPARh1eg9zah6ii+cQhQpGFa2348HzDYUBxKlAvofnEZCRM
iaYr2kMCMzKaJKC8hlue7Q5HaTCk8kTG/G1OBuYrLFWVra7RYkJV3vbqwKgdWdsC1ET++6OyxKCCVpYUHL5tu8W+v893AwXKS2So7mgMfcf7ZigYx3D/J/uOoduvkkLO
imwCyuUgSJzdNdWn1mcBysN4xfXnrZS8v/num2K0qNi3mSSfLSARcoabbMIjOJDfBtvHXOaTNohnt2G43uJ5PX79xoo/6Qu195827gVBf+9uFy7txBzP6Zz2XZgCnNFm
YGq27kuNRTfOQztvyjeD2hgR2xXDyc35v/+x3abIb4izkeUJMNYnrFx+zzHkakhPxrqlDRFDM4VekkAFoPghdfZfq07MApPCfLxbhk/JS4c3f14fFH86/w2cL48aDYhG
w0CTrRm7EZ1/uWt4Ud2LmgQXNRJdDsI9PRff1EYe41I7OZi0BvupsnSJD1tPQjjuMSGjcjWH3vGcxryv6it/wzHElrClgAoVM6rmRLT92tf5H18vvwqVg3IKV5ivs3ik
H+sVmvMKpNAEfnrB7Z7CGdOwCao95KeCi/nOQHhnkzZUv27LvQUL1c/ntTmWogj1PFXdVbtxFepJZP66g/nVKqnKl12w3/RkWXbG2HzrJSBNe7skDS+Q6kbld1qfr3tO
z9zKHfERRpo5MxNsYvilWmXzZSXzHNbq/yAGJlujqjfCbQcwVUWNURxkzPOQpG3pxb6/z3cDBcpLZKjuaAx9x/tmKBjHcP8n+46h26+SQs6KbALK5SBInN011afWZwHK
w3jF9eetlLy/+e6bYrSo2M22rMgUCc289S+rtcgOJj4feKkOC+6sSX6kuyc2oQ0HxMKI8pDTsHTAAYa9Ry7am4QvsggK03c3rXUqxEd9Ru/KFBhS4kozqPVJbtX6uyT6
yrWl1Yc9jvzkoebAsNT8DpyZ8ZoCi2j7WXFQYBYwcoizpcMzmhOQTlp5GiRJnwNYqHXx4aVIhWBF1HKVz5BPepyZ8ZoCi2j7WXFQYBYwcohtT/cC3ccdSgmz/dVhCTW8
l+qVjvEZKiHKj3AwZ0nNHJyZ8ZoCi2j7WXFQYBYwcoib7pwvMgh34M4qNN1aV4y2e2c9y9IPLAMn3GFUo6HDxT1oTPaT2lxds+LyD42iUDfail28E99+wg/W/uK2yLR8
MmF37jlK3AnpO4WymR0ZWRTAUdExGH+mDKIGbzdggHZdvXPLMV0cw0du8YzldjwuNnlzPq/hK6t6UeqBEASytFzWMBSgOoE6gSOCmFUqm4q86f8O7htU2jHKhyAfoRdF
MZriW6sBHaZY3e0W2XFKb8a6pQ0RQzOFXpJABaD4IXX2X6tOzAKTwny8W4ZPyUuHN39eHxR/Ov8NnC+PGg2IRsNAk60ZuxGdf7lreFHdi5qF0vC0cGkYnJcY7Z6I+AHI
jGfoYGVDhkskHfFPMYqGgMkcOIm0U0hekOiAW4PkZrCu6/LIxH9svswcTn1m9sWBUn88uuBDEtPJJ+s6Vy3SJV29c8sxXRzDR27xjOV2PC42eXM+r+Erq3pR6oEQBLK0
wqPw5CJLYUWWRKkmzXhu70S0oympk2Wb3M4OK656laldvXPLMV0cw0du8YzldjwuNnlzPq/hK6t6UeqBEASytA29mxthVMiEhjOqpSfw3h8XWo8QOn3yJfaJqQXCtVmB
Xb1zyzFdHMNHbvGM5XY8LjZ5cz6v4SurelHqgRAEsrSCAqaMDQrNHhXwtG3vxw70UIYHoLjhxJV/r1J9FeQa8fzwxB6sVPMLyLOaYqfxm3Oze6G5LTlpIP6cwQ9HIOPV
xYZICqBGtB6VVnOsjp6s7ndE48XHt7GBrIzJf1GPtsAtGw0PCF1cAUm1C+9L4u3Kf3ljlEZ9JR6b9dEMg2aqJS/MNzMfl0c8z7+hsIbrXExqsWAJuVmyGvUmGaDgwQK0
s3uhuS05aSD+nMEPRyDj1cWGSAqgRrQelVZzrI6erO53ROPFx7exgayMyX9Rj7bALRsNDwhdXAFJtQvvS+LtynEHFErppmd2Lz2lv+fbEYj1afC3N9kGF7REmQ1xsxQU
IIv4hZpCZXviI5crqhlXrcw2+0CToRJCsvlWhn5N8vlZAQsW/mfx/ZM248LaiUvIhLFEsuSi05pIZzxqztlf8dL0NyUqqmPT+HEKPWivr2lblcCZSh7LxlHXnPc4CfPj
L3Qz9X1IPj0mbUa8TXAGKtOMIQSnCHoVvPwtGDRvghr3KNeETLzgcnQ7fcZT3ljxWQELFv5n8f2TNuPC2olLyISxRLLkotOaSGc8as7ZX/HS9DclKqpj0/hxCj1or69p
W5XAmUoey8ZR15z3OAnz4y90M/V9SD49Jm1GvE1wBiqlxteewgOt50vrWtJON1xt9JOmEDXyoQIKUfzB1GqTeh94qQ4L7qxJfqS7JzahDQfEwojykNOwdMABhr1HLtqb
hC+yCArTdzetdSrER31G78oUGFLiSjOo9Ulu1fq7JPodYJjhjAwEN7EJgU2DTt+9WfS5sFGfRMDZCGlKeqjj2USQIG1JUAE7jlHwvtN6vhpjfT7Okme8IvOUQmioZFDO
8ZkcHRIwyQSIyTLThunP3QD8MimiUKzmAFmkik321+KJ7LLf7XXqHv8pMJ1Qc384yCG71MOOtc2dTsG0UYHmIz+weKxefITRZ5UuIugH0J1debuWM9GQT0QV5SXpFY0X
myPpjN/jiMUqpJTIbvM42zTLKHT9tINDpIOhV1mZjftJpOzMj/yzR+sp0xnL8Li+q3Sa47bTrGgA4mOjOT3Rr003QcZd1UsoZo4oBoaE6n70nhfLLzWBKbGMeAKCpAMO
rSxJCmdo4Vy5G8ZU+jb5FR7XiDUZgfSHix9bLxm2wVkYHvsf5GLe0t2edTuvwkJvwTOsN6Xr9drrzMJgB3ARtQA4oF8WTFAw2FeaIuQNFZH5aJitZZ8o9FrOQT6VKvJF
us47RsEwUX1D51MVb8t1Ksgyj2YeOPlcohDVFnTNT/24DG3BLdwdNEvA0vspgS2rgpuwEt34Z8r97z20GbuppnP0AX8uLNZ+9N1KpgVY9QbjoY62Wru0MBPPXYJzG6Xh
ZigP9/FrkP+qa5izOBahgsghu9TDjrXNnU7BtFGB5iNFgB06EEVMhLZrMy01CrocIIv4hZpCZXviI5crqhlXrR4YpCoQjbLbPWoxKzJo+Z0TL6tf04NPgH+vCaoAdQTq
A1UdnG9Q4Sl8nnHOS5G76gsqtOJAG83XnHPKembSHIlVzdpDUs5dM96giH+z6uI/T471iFw7YcwrtrPjsRZuxMghu9TDjrXNnU7BtFGB5iN5MLGLvbiECao1V4LO+xtf
yo9uQlUUmiECJbyckZKUiawRckptv6ma2gtKIe0mcuP7j0PBEMk2P8v9GizxMvkFtvniBMMegANO3ptBGO6ohtId7QG1ElGE5vvkz/Tosf3A6iGQIk9/K4AHE1BnZ2s7
M6k0fanmHuoru0iCY98wQ+x+vvSywjES9kpc+s6FhLRfPIm4RJiGU6hlgG25jFkvSStZ4bEk6M4R1VAKsSWEq2SSdsCJg74/R7snMXOwc71F87NlWpGJK1MFDB8YDx0H
YMVkmuWPMb5IONJjrCIqLzhHTkxhcKFCsePvAI6Q1Lt5PSpTr6cmqu/g7fFTpy8BcdOwFk9lnsWLsL3/muCqVMPv5T95EcJNAPHCG12y/Zjdgt6wCU4j3I5PVnb2pbo5
2vbtj65XEsDGi305XpA7D8wWgUMXWTVzY97zTlc60K0Ix6Ve5jYJr8ORTQuvh+hwGZfpQv2Q80ojIziSg8o0U1hRXrGB5LRsR2KRIureqPQrpYfSX1L5P3i8LHFTZP22
U68r3JcRmYkg+L2BDBKdVF7yKW9i+F07HSgTgxQFAHIyN/mJb13oaQMfLt9bHhnzG08JHD87nW89oL8CdhdD1BXJadX1ib3i6mni8t3+mUb6xvxcaHosKZTOSsOU1QwO
nIYn2ZMgVuSHfjeWXIKfdHdoQGY4lnfXs7KOmoBw3wr1r2jgLRVNS/HqA+r3l+YfhMd3qtW5XDgZXNk5rl6RRrZPfAtN9GTdZucp8rIl/AO3l36g0qrlqQEQsAGQx/uH
7LYctKoMc6k7jKklhcUE2IyBChyLrx5jmXws+GvkzyIDTqrjwfHBNqw0NPF9HICgHBKf3XvvI1QmVPkbEThDwnE2ZOjPKs+cmcw9gmJ5eYV0tF/Ml8q+Uv49uVBIFQG1
l7zuVQf4HT1id9hnfAhuAcgyj2YeOPlcohDVFnTNT/0lbbbhsbm0slngRKvARnqPfGGJJGbIA+2xs5fFqdQ/o6vHZrXHUPSodvVQZPy3wANSY+3c3neQTqQ2BOnRi51y
AgmDleCXxtCBGrUwBGQ8RuIZXFj+TM0g/yG8bpDqs2tTJiPI94niD6nVzmGh6yFD1EZmFD40ajXoRQDlIbzO5pMvgddD/CW+rSnB7XtQhnM7oeBURpzihLXJC+iSlM7a
qq9GUxASCTTOmP3K1jhM0Ssc643vxecFNSfRtb2b3V8r25FgHUwak/Y52YK/nCVYmXQZ6PSEdauWjNsWGLN6yymNWX/36R7gfrdxy3vFHixh7m9hW6kGuklFOZWKy5DH
WQELFv5n8f2TNuPC2olLyISxRLLkotOaSGc8as7ZX/HS9DclKqpj0/hxCj1or69pW5XAmUoey8ZR15z3OAnz4y90M/V9SD49Jm1GvE1wBir1nKTDpGfRTLKpVbIY0d+W
BqNtSSmMDBJiwKY0/NaMClWE7PBI6EPgdmjKhDnu+QXtPmimPWeFyuR7CoDvDg/RJPsTqUddPqzMmwInI1A2UrN7obktOWkg/pzBD0cg49XFhkgKoEa0HpVWc6yOnqzu
d0Tjxce3sYGsjMl/UY+2wC0bDQ8IXVwBSbUL70vi7coY68H5x1OFMI38+2cAvqUL4buRwVhLdfLrgVnZx9I2k6IMV5MZSbPanZ/0qh1PPhi2R9jUsmX/W6UCBWyqWI2J
IhP2P0ZGkAbQ8THOQc4K4qQtlgvq5Hp/YwOX8NE5+nnrx9HBQiSZCmL4VWEP1fsUPFXdVbtxFepJZP66g/nVKqnKl12w3/RkWXbG2HzrJSBNe7skDS+Q6kbld1qfr3tO
z9zKHfERRpo5MxNsYvilWsukrewpxK97OhV9/mvf4zVc87IOTcgLSaToZt+lYHjUPjgeYGg75D6NgYgTLYWWwm1PVG/eQM1Mts3i33GohtocU+VhbTgQOcJjFYnuFYzH
75hDSmaNh1GI59Ls6CRU4Po/zYjUtGdAJihn+lK0LjwpSCHXzB+SRXhODlnT4VF17EXOGu/j8vMenfeI3AE0TsROWIPqqK6nnXL4mrsDCJP+qwN3BzD96QwImyy37IBk
rggwLrGV2pVqBHbWejMPZOi/hO5WbRVRyCXSLysoNgqf1b4ms4jHm2DlgudsQFsNZ9mVT7SVRohCNCuzwokqwvTe28VwLA7Gr1iZUbyT1zByn0EB7W1neic2RU7pUpJb
qT4fCpsUiI125SFiSA0PNq3F75sspHOCwJ64J6v6T1LjwsvAit7u+kuRabzahUnjwCwlJ5DiHDS9a1EBad3hiycrg+FUB/V6J3bc+ICS+YedG77qT0pL/25BPXQ9DqBy
zmhHYjYrWLLO5EHpZPREXle+tmmI8OY5Iny2Uz5HhRdsnytP8jJBpGPUPdY4cmvEBTu1x3wlS+alZjpjAjiesST7E6lHXT6szJsCJyNQNlKze6G5LTlpIP6cwQ9HIOPV
xYZICqBGtB6VVnOsjp6s7ndE48XHt7GBrIzJf1GPtsAtGw0PCF1cAUm1C+9L4u3Kq1GOXK65ahbU07tsTrf2Psa6pQ0RQzOFXpJABaD4IXX2X6tOzAKTwny8W4ZPyUuH
N39eHxR/Ov8NnC+PGg2IRk9YYv+PPqJiOSM+Wl5gqVBptieiqqLJ4tCYKHX6Rno0WXQVwrPHT/yd6EbO1LN1X7+plDmE8EQz/nEY9rk/gbn36CkqBLVwG89HUkKjc+4A
jqON4P+jJtle6sXdARQTE/tQfx02f8/IPBfmkDiknVCUXxDj1sgNV2SZvRrDpvPDLI8P43P0uM/NdAfVXFREUYJ6kqfY2ARnLuZi6XU57mD48HzDYUBxKlAvofnEZCRM
iaYr2kMCMzKaJKC8hlue7Q5HaTCk8kTG/G1OBuYrLFVUs/262kiC9e4jcFnQENLt1IHMg1bw8M47SJKpBpC1qSE0AS7WJOaQ0RqwrafqV6/bCIT747TZSvjvMWbVJB4S
kuuhhq4mVW1kDGh6tUBNxyGm6FinxMvWYzd1Xu10V2vK77RB6IEtqVOQ2ENBHstx59qk97G2l1H47CzM1D1BWlgF9GkqvI3T532KH4N1qB3FDAtjstydgkH9WkIZMYIi
ms6HN3nXMcCrWnmM2pYlZH5g3B7IqptlP6eQom2zXTx0DQ4txMGz/3HQLI1gnwMlOz4VyjAcg9Zlj+cwFwFDXrx8oZcO/gnv7M80supvdcwAPM4tEjK7iYsN5uMLgI38
U2lYzf74CGZmoaFRFGl6ILvhaScnS76hKDNCiqUpDRPO0rq/D5zDIfJsFQ3sO1YDTNqqeiZITbjceBEELp//w35g3B7IqptlP6eQom2zXTzjtT4V+9ZWmf8t72jDAUvA
ZOfDb0YOZlyjO4u7mVZnNvO5YvHEvGP/yqh41g/Z9kWb2BNh55TQk+b8gwIF7NFpMcDcrS/rGEq01gip2YmxVr1kVCqlYRYZC07/5l5IFE4rRQPV9SFNuPBfOqrVkV3m
P1gDmwJmD1qmgbe1YadBdapStNyb72EsrtPz09QI5ErLNh5L7cQKkjS8IhE2+A8nLq+mLjyMDe+bNcrJvnp3IZt+SYUIxU2zCShKWGPoEChwIB/84iOtkDuRBUr6IV3w
iY1Onv3JhWzY+O4XzF4dg/9nKzqRzw+XxL75ltoOZbnHLMJmii5i8NmeuMHFBGneImRQODrDzM/sLi+UPFilQ+nLUZOXAuwW0BNj65bQxZwSbP0aBPHHUt8wvmS97itB
+X5Q8pmLQHmBbvk7WupHf/X438VFOgyYMQ8w6MjxT1Coeva8QmGqmV/J64gY0ZpX1jnBuTKmRns7OgZQOPqQAwlmeBa6eocWFRqHMLz8F1l8pIVDRagIAplVl/6g4xSv
yzYeS+3ECpI0vCIRNvgPJ1m25zGiYl5VhjD9X2DefC8Swq/FXEc10MuX+KMqCXsY8Wqh92/Dvq0tmiwRPzvENuYCAH2cTccs3aHvhiTPe9R1yfulOp3DA2prRUHnM6AB
m7OUpyqr9qjffPe27Ox6Aui5hxjxM5N2z5cQdnIJBi3FRA6D96LuQTVMZEqNo/PxQ8TmkzC3Bj1ixAx3wnt3qCmfZ5sNkYGfmJxTfC5nSPu54mUrNogou2XnrEaCECRU
m7OUpyqr9qjffPe27Ox6ApQHQaYbbvQf1Pt9avxEeOwqHDYBrYd4vbqJhccE7sMpol9b4BpyvukZDRA5O59XK9h9DEmmf8SwWgh0ZB0+gLD1ylHAa9zNQQ54aMqZQ7Te
JGxTZSak945RYVqXm/ZZMwfYHjb9cFZ02+ldvTQS4SiWpz3iY67U8zx5XBJSQO2umJJA/611Sddj53Zc5IDdmpzP04XSkbIjZF796FAq/6jObm40/VEc4tQ6W/+I9hVQ
4NxvQX4dX6TvlL9w5HXwf3dGaucvJSUEa8kYv5OOGG06hwS3MdyRcT/8X5kMdS10yogm0Sa9h4GMq195YwJtiCbaj3E0QhDi37c8qTt2pJKuHi1w8/uOCcDGu+LNo49D
9eG2OLGIKwH00Q5QBYbs4JoiPd+tizCzzWWfZtpSw0aaIj3frYsws81ln2baUsNGCBzMADeMeWn4Jr2PCFcDIpuzlKcqq/ao33z3tuzsegL3rUqOOiTSIdhTIMg5HViu
w5KLT9SFoznQGp/mk7winyfoJ/CXL/mF5JwPsuxnmLTRWk8HZ9TQ95vgPDt7XVl1DvotatZigs4bDxWBgEKgXxnNz7LcM1Phn40OlxkidLaHSeHErXIDOUTwQIYowV6B
hLvQEQLaeVmfrExn+Dr+3MkIle3xS+tpolmWjghZocNOo9QUB4hmFuJ02MInEhWc4XjxK32l1WL6V7sqPmWZ+TNSCOSt51kl2Cl8h/O2snTRdGxfbWaY8K/Ao9y1gs3c
rAMuIFCArwe5VuXT2hX7NS6SQX7zUY+yfrFiRq75Bf0RlkG+x7k2y4Nf+H67/0WfaRA7pmL3TRA0PXPayCQra1prkOP6vRsYDREA5wCq9G7/rcHltj5Xc7kPP3FiI8eS
iqufVS6TOUhCNpjOJbgnTm6KrJlHhzbSxI+D1/Q2fd73IKyql7f7oKt/zgXwYEL8JUchTzuuZdzmhYdC/uc4Wj1QEBICPyf8egYy8/qqHPPs6dcM2krk4xy9ofvBdlZt
ix4uDubYCxHC2GXdOXHmkBnVB0V4f17dBuBdSYzRb68CxfnE0AiPyGpIn3/t7QfYsZz40R6ZEtGPW51Tk8A+8MMpt/Vo7UKrswexZSU4pLKLUW/QwZm+IXEBpzcMZEP2
Sa9jsqCj+0kuJ6lw8ejcTbX8DFl24T99tEYbRF3hrx9kVpRd6aoDH8nXdyfrOWx1+zqC3u7kmfui84FrM34lanteYyhrLI+C5J8UDDx2D6/aX5eRXQhhP63yHkSVXBkD
xbvgwn/Dn7RF9hhkpSFAAdZ2PS8H36DETzePr5Q/YLk3E/6LBchmsRX2/fYXTVBhUzunwoiEbupzfjAxoFQgarxGRurpa6xbNvFnJDsJfTEPIZLNt032S30Rxa2yU7gH
BqIhCfexYwcDEz5wt/9b1xrbJvFYqFamSHjoEzCZxJqf7G1kmbXYD1/Hwf801xve+6w6dSlSm6Kr4rbJD4GzSE5VV/BUqdCHw19+i6ILooQ1yYl9EssN1ahYxH+flUqz
QtPn5+TbV4Zvkn79E4hAAwGlnsRRHhwVn2nz1vHqhirCSqQdK6eASRlcfAEYhroKqp6cXVbtA6A2QjeYwFyCsai+JN7IsyVtG9dggvy8rM3U2yXvi8HZYuIE283f2mJZ
JxUfKCQlIaqfw5V006IkZ41zBPkTFGYnSjYIz10ya1D4ddrb/VnYU791mN43qiReyR6DFYwVcm0Xjwlua8sm0CPNI5/NJx0LXaJLd+SyjUJdPl6rStOxCLNwHpFwjOrk
TAjTA/mH7hb91fJ6eUMXGZxmHqoafC3FVXUf3N9EtQyfiUZg4+nlg9SxG86P7FbWJcvX5l2sw+HUaLwBkIn8EYSuvt3MhFZMu1ODfWZeUgtnupMOKb8bh88ywZI5hEWI
JcvX5l2sw+HUaLwBkIn8EUP5pBo3ddFBTMFnnI67A1k8BN0uqCsZaO4xnML2SftP+bNs61L5B9dlMnmDVUPMbl3jtC1P/IZi6a02WQux5pkHyVFkGh4GxZmJM7psuNwy
rS0GmpsCk6T/xZ0WT5x2cA6YWSkRynBI9i5EiBDC3FFlUsMBwB+DqxgJGGOcwS6sjuJfKqjw5j+FjhmMd1XleqOrT4d0nMTC+O4riyUyG+VST8V24SoDc83i+GeKwaDe
HHD9VYQGZm8xQyQ8hwerh50xZpjkZIiBukIG2bAhiebnwojcwcKPYkZ9uHqsuacwDQ4RhvJRb9lJAdC3gGwTubkey5LxBNm24toVlkYpQErE4AWZXJiIaxNp6ZktBHnD
qIEkOH26tSb3deh80LsNUDo7X4f5uHU9RO+rrDEq5D6Ad0veuv3qbA2emRxHB281NNCTFJQYt8o0IWti/DNiVwQRuXsXVcNuNwF8171OU+zawhr7z602iNQMdyJI+I7p
aoHBG7OyUsV9iWABA+O7lt4DGngfKKoOAdlaAOO2C9/1B6JO4HNKijJ/Hr7AXcaTxOAFmVyYiGsTaemZLQR5w36ROTa1ev9YWXY91+oDCH3UlKD/Ut5EwQqUwcvKhS+4
U+4mUPNKbJxFam7p+QPKY5/HfAtwGn6C07s5+Bzu6zfpv1SKFXc/643bAW2JiXtN0TooCBZYm9AePULi8dyT9DIWEOOAduf4QZ3aZ/DeuaOZP5TyzUH/LBKtcaOSgTK6
B+Z1Si0vwBV/Ffq8t4z565WJAgxUu1EV1mJSML89TXSeE0vuhLm49DVYu5AGZu4LB+Z1Si0vwBV/Ffq8t4z56+q/Vcsu4DF01xG/u8Qt0R88g/824FPy3yW0dFq36xSi
dwCGjPIjEsxbumHmKEXBfAioNL4LpRu4qsmXBwhOIimKZcfClFqTpJzAaxmni4S7gYW5MKk5YfCHX8yESBWPlpVApCgkf4Tmb0z9VpiLGGyr8JinN9xZcYadpXQ2dhth
LFIzBRkvE72jYLtVIwD/va2hQtrFVEiiCzCCFaeBZT+3rGVBtkbAvPjMDJdZFyLbflYTx8TIrwItNFHXEieNLWp506MvCkkn9jCfwIfI8D6vNo0IPqAyCIUCiZmPLydt
fAGxopsBcL7c4aIPml8uGukjzHqalmxxcGC+R9/RFjPhsgeBRaLW5blz0nv6+daopkH23IDqfDxo1P9GUU0mAlBpJzGHlYF3RUl6WC7nDCz/jVE0y2cb4JMkr8GrEu5+
k/lRw8+3lXtHdI1XT0c6Pd8nhvFhBmBUmqe7sEsOVZhST8V24SoDc83i+GeKwaDeLFIzBRkvE72jYLtVIwD/vVzNHBDpKSAfMWqVo6ZY3m0nyQ5p7SzY5X5Kjt89xOtV
lL9FQN8JRK1Gab1GxmusRQXznXbX2gAL8VuoJ95F1YP2VoWL3frBdGNLwRJDLAw8
`pragma protect end_protected



