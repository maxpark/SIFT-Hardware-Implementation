`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:34:16 06/13/2022 
// Design Name: 
// Module Name:    dir34_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module dir34_2
(
    input   [7:0]       a,  // Addr.
	output  reg [4:0]	spo // Data.
);
	
	always @(*) begin
		case (a)
			000: spo = 5'h1b;
            001: spo = 5'h1c;
            002: spo = 5'h1d;
            003: spo = 5'h1e;
            004: spo = 5'h1f;
            005: spo = 5'h0;
            006: spo = 5'h1;
            007: spo = 5'h2;
            008: spo = 5'h3;
            009: spo = 5'h4;
            010: spo = 5'h5;
            011: spo = 5'h6;
            012: spo = 5'h6;
            013: spo = 5'h7;
            014: spo = 5'h8;
            015: spo = 5'h9;
            016: spo = 5'h1b;
            017: spo = 5'h1c;
            018: spo = 5'h1d;
            019: spo = 5'h1e;
            020: spo = 5'h1f;
            021: spo = 5'h0;
            022: spo = 5'h1;
            023: spo = 5'h1;
            024: spo = 5'h2;
            025: spo = 5'h3;
            026: spo = 5'h4;
            027: spo = 5'h5;
            028: spo = 5'h6;
            029: spo = 5'h7;
            030: spo = 5'h8;
            031: spo = 5'h9;
            032: spo = 5'h1b;
            033: spo = 5'h1b;
            034: spo = 5'h1c;
            035: spo = 5'h1d;
            036: spo = 5'h1e;
            037: spo = 5'h1f;
            038: spo = 5'h0;
            039: spo = 5'h1;
            040: spo = 5'h2;
            041: spo = 5'h3;
            042: spo = 5'h4;
            043: spo = 5'h5;
            044: spo = 5'h6;
            045: spo = 5'h7;
            046: spo = 5'h8;
            047: spo = 5'h9;
            048: spo = 5'h1a;
            049: spo = 5'h1b;
            050: spo = 5'h1c;
            051: spo = 5'h1d;
            052: spo = 5'h1e;
            053: spo = 5'h1f;
            054: spo = 5'h0;
            055: spo = 5'h1;
            056: spo = 5'h2;
            057: spo = 5'h3;
            058: spo = 5'h4;
            059: spo = 5'h5;
            060: spo = 5'h5;
            061: spo = 5'h6;
            062: spo = 5'h7;
            063: spo = 5'h8;
            064: spo = 5'h1a;
            065: spo = 5'h1b;
            066: spo = 5'h1c;
            067: spo = 5'h1d;
            068: spo = 5'h1e;
            069: spo = 5'h1f;
            070: spo = 5'h1f;
            071: spo = 5'h0;
            072: spo = 5'h1;
            073: spo = 5'h2;
            074: spo = 5'h3;
            075: spo = 5'h4;
            076: spo = 5'h5;
            077: spo = 5'h6;
            078: spo = 5'h7;
            079: spo = 5'h8;
            080: spo = 5'h1a;
            081: spo = 5'h1a;
            082: spo = 5'h1b;
            083: spo = 5'h1c;
            084: spo = 5'h1d;
            085: spo = 5'h1e;
            086: spo = 5'h1f;
            087: spo = 5'h0;
            088: spo = 5'h1;
            089: spo = 5'h2;
            090: spo = 5'h3;
            091: spo = 5'h4;
            092: spo = 5'h5;
            093: spo = 5'h6;
            094: spo = 5'h7;
            095: spo = 5'h8;
            096: spo = 5'h19;
            097: spo = 5'h1a;
            098: spo = 5'h1b;
            099: spo = 5'h1c;
            100: spo = 5'h1d;
            101: spo = 5'h1e;
            102: spo = 5'h1f;
            103: spo = 5'h0;
            104: spo = 5'h1;
            105: spo = 5'h2;
            106: spo = 5'h3;
            107: spo = 5'h4;
            108: spo = 5'h4;
            109: spo = 5'h5;
            110: spo = 5'h6;
            111: spo = 5'h7;
            112: spo = 5'h19;
            113: spo = 5'h1a;
            114: spo = 5'h1b;
            115: spo = 5'h1c;
            116: spo = 5'h1d;
            117: spo = 5'h1e;
            118: spo = 5'h1e;
            119: spo = 5'h1f;
            120: spo = 5'h0;
            121: spo = 5'h1;
            122: spo = 5'h2;
            123: spo = 5'h3;
            124: spo = 5'h4;
            125: spo = 5'h5;
            126: spo = 5'h6;
            127: spo = 5'h7;
            128: spo = 5'h18;
            129: spo = 5'h19;
            130: spo = 5'h1a;
            131: spo = 5'h1b;
            132: spo = 5'h1c;
            133: spo = 5'h1d;
            134: spo = 5'h1e;
            135: spo = 5'h1f;
            136: spo = 5'h0;
            137: spo = 5'h1;
            138: spo = 5'h2;
            139: spo = 5'h3;
            140: spo = 5'h4;
            141: spo = 5'h5;
            142: spo = 5'h6;
            143: spo = 5'h7;
            144: spo = 5'h18;
            145: spo = 5'h19;
            146: spo = 5'h1a;
            147: spo = 5'h1b;
            148: spo = 5'h1c;
            149: spo = 5'h1d;
            150: spo = 5'h1e;
            151: spo = 5'h1f;
            152: spo = 5'h0;
            153: spo = 5'h1;
            154: spo = 5'h2;
            155: spo = 5'h2;
            156: spo = 5'h3;
            157: spo = 5'h4;
            158: spo = 5'h5;
            159: spo = 5'h6;
            160: spo = 5'h18;
            161: spo = 5'h19;
            162: spo = 5'h1a;
            163: spo = 5'h1b;
            164: spo = 5'h1c;
            165: spo = 5'h1c;
            166: spo = 5'h1d;
            167: spo = 5'h1e;
            168: spo = 5'h1f;
            169: spo = 5'h0;
            170: spo = 5'h1;
            171: spo = 5'h2;
            172: spo = 5'h3;
            173: spo = 5'h4;
            174: spo = 5'h5;
            175: spo = 5'h6;
            176: spo = 5'h17;
            177: spo = 5'h18;
            178: spo = 5'h19;
            179: spo = 5'h1a;
            180: spo = 5'h1b;
            181: spo = 5'h1c;
            182: spo = 5'h1d;
            183: spo = 5'h1e;
            184: spo = 5'h1f;
            185: spo = 5'h0;
            186: spo = 5'h1;
            187: spo = 5'h2;
            188: spo = 5'h3;
            189: spo = 5'h4;
            190: spo = 5'h5;
            191: spo = 5'h6;
            192: spo = 5'h17;
            193: spo = 5'h18;
            194: spo = 5'h19;
            195: spo = 5'h1a;
            196: spo = 5'h1b;
            197: spo = 5'h1c;
            198: spo = 5'h1d;
            199: spo = 5'h1e;
            200: spo = 5'h1f;
            201: spo = 5'h0;
            202: spo = 5'h1;
            203: spo = 5'h1;
            204: spo = 5'h2;
            205: spo = 5'h3;
            206: spo = 5'h4;
            207: spo = 5'h5;
            208: spo = 5'h17;
            209: spo = 5'h18;
            210: spo = 5'h19;
            211: spo = 5'h1a;
            212: spo = 5'h1b;
            213: spo = 5'h1b;
            214: spo = 5'h1c;
            215: spo = 5'h1d;
            216: spo = 5'h1e;
            217: spo = 5'h1f;
            218: spo = 5'h0;
            219: spo = 5'h1;
            220: spo = 5'h2;
            221: spo = 5'h3;
            222: spo = 5'h4;
            223: spo = 5'h5;
            224: spo = 5'h16;
            225: spo = 5'h17;
            226: spo = 5'h18;
            227: spo = 5'h19;
            228: spo = 5'h1a;
            229: spo = 5'h1b;
            230: spo = 5'h1c;
            231: spo = 5'h1d;
            232: spo = 5'h1e;
            233: spo = 5'h1f;
            234: spo = 5'h0;
            235: spo = 5'h1;
            236: spo = 5'h2;
            237: spo = 5'h3;
            238: spo = 5'h4;
            239: spo = 5'h5;
            240: spo = 5'h16;
            241: spo = 5'h17;
            242: spo = 5'h18;
            243: spo = 5'h19;
            244: spo = 5'h1a;
            245: spo = 5'h1b;
            246: spo = 5'h1c;
            247: spo = 5'h1d;
            248: spo = 5'h1e;
            249: spo = 5'h1f;
            250: spo = 5'h1f;
            251: spo = 5'h0;
            252: spo = 5'h1;
            253: spo = 5'h2;
            254: spo = 5'h3;
            255: spo = 5'h4;
            default: spo = 5'h0;
		endcase
	end
endmodule