`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:34:16 06/13/2022 
// Design Name: 
// Module Name:    dir28_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module dir28_1
(
    input   [7:0]       a,  // Addr.
	output  reg [4:0]	spo // Data.
);
	
	always @(*) begin
		case (a)
			000: spo = 5'h17;
            001: spo = 5'h18;
            002: spo = 5'h19;
            003: spo = 5'h1a;
            004: spo = 5'h1b;
            005: spo = 5'h1c;
            006: spo = 5'h1d;
            007: spo = 5'h1e;
            008: spo = 5'h1f;
            009: spo = 5'h0;
            010: spo = 5'h1;
            011: spo = 5'h2;
            012: spo = 5'h3;
            013: spo = 5'h4;
            014: spo = 5'h5;
            015: spo = 5'h6;
            016: spo = 5'h17;
            017: spo = 5'h18;
            018: spo = 5'h19;
            019: spo = 5'h1a;
            020: spo = 5'h1b;
            021: spo = 5'h1c;
            022: spo = 5'h1d;
            023: spo = 5'h1e;
            024: spo = 5'h1f;
            025: spo = 5'h0;
            026: spo = 5'h1;
            027: spo = 5'h2;
            028: spo = 5'h3;
            029: spo = 5'h4;
            030: spo = 5'h5;
            031: spo = 5'h6;
            032: spo = 5'h17;
            033: spo = 5'h18;
            034: spo = 5'h19;
            035: spo = 5'h1a;
            036: spo = 5'h1b;
            037: spo = 5'h1c;
            038: spo = 5'h1d;
            039: spo = 5'h1e;
            040: spo = 5'h1f;
            041: spo = 5'h0;
            042: spo = 5'h1;
            043: spo = 5'h2;
            044: spo = 5'h3;
            045: spo = 5'h4;
            046: spo = 5'h5;
            047: spo = 5'h6;
            048: spo = 5'h17;
            049: spo = 5'h18;
            050: spo = 5'h19;
            051: spo = 5'h1a;
            052: spo = 5'h1b;
            053: spo = 5'h1c;
            054: spo = 5'h1d;
            055: spo = 5'h1e;
            056: spo = 5'h1f;
            057: spo = 5'h0;
            058: spo = 5'h1;
            059: spo = 5'h2;
            060: spo = 5'h3;
            061: spo = 5'h4;
            062: spo = 5'h5;
            063: spo = 5'h6;
            064: spo = 5'h17;
            065: spo = 5'h18;
            066: spo = 5'h19;
            067: spo = 5'h1a;
            068: spo = 5'h1b;
            069: spo = 5'h1c;
            070: spo = 5'h1d;
            071: spo = 5'h1e;
            072: spo = 5'h1f;
            073: spo = 5'h0;
            074: spo = 5'h1;
            075: spo = 5'h2;
            076: spo = 5'h3;
            077: spo = 5'h4;
            078: spo = 5'h5;
            079: spo = 5'h6;
            080: spo = 5'h18;
            081: spo = 5'h19;
            082: spo = 5'h1a;
            083: spo = 5'h1b;
            084: spo = 5'h1c;
            085: spo = 5'h1d;
            086: spo = 5'h1e;
            087: spo = 5'h1e;
            088: spo = 5'h1f;
            089: spo = 5'h0;
            090: spo = 5'h1;
            091: spo = 5'h2;
            092: spo = 5'h3;
            093: spo = 5'h4;
            094: spo = 5'h5;
            095: spo = 5'h6;
            096: spo = 5'h18;
            097: spo = 5'h19;
            098: spo = 5'h1a;
            099: spo = 5'h1b;
            100: spo = 5'h1c;
            101: spo = 5'h1d;
            102: spo = 5'h1e;
            103: spo = 5'h1f;
            104: spo = 5'h0;
            105: spo = 5'h1;
            106: spo = 5'h2;
            107: spo = 5'h3;
            108: spo = 5'h4;
            109: spo = 5'h5;
            110: spo = 5'h6;
            111: spo = 5'h7;
            112: spo = 5'h18;
            113: spo = 5'h19;
            114: spo = 5'h1a;
            115: spo = 5'h1b;
            116: spo = 5'h1c;
            117: spo = 5'h1d;
            118: spo = 5'h1e;
            119: spo = 5'h1f;
            120: spo = 5'h0;
            121: spo = 5'h1;
            122: spo = 5'h2;
            123: spo = 5'h3;
            124: spo = 5'h4;
            125: spo = 5'h5;
            126: spo = 5'h6;
            127: spo = 5'h7;
            128: spo = 5'h18;
            129: spo = 5'h19;
            130: spo = 5'h1a;
            131: spo = 5'h1b;
            132: spo = 5'h1c;
            133: spo = 5'h1d;
            134: spo = 5'h1e;
            135: spo = 5'h1f;
            136: spo = 5'h0;
            137: spo = 5'h1;
            138: spo = 5'h2;
            139: spo = 5'h3;
            140: spo = 5'h4;
            141: spo = 5'h5;
            142: spo = 5'h6;
            143: spo = 5'h7;
            144: spo = 5'h18;
            145: spo = 5'h19;
            146: spo = 5'h1a;
            147: spo = 5'h1b;
            148: spo = 5'h1c;
            149: spo = 5'h1d;
            150: spo = 5'h1e;
            151: spo = 5'h1f;
            152: spo = 5'h0;
            153: spo = 5'h1;
            154: spo = 5'h2;
            155: spo = 5'h3;
            156: spo = 5'h4;
            157: spo = 5'h5;
            158: spo = 5'h6;
            159: spo = 5'h7;
            160: spo = 5'h18;
            161: spo = 5'h19;
            162: spo = 5'h1a;
            163: spo = 5'h1b;
            164: spo = 5'h1c;
            165: spo = 5'h1d;
            166: spo = 5'h1e;
            167: spo = 5'h1f;
            168: spo = 5'h0;
            169: spo = 5'h1;
            170: spo = 5'h2;
            171: spo = 5'h3;
            172: spo = 5'h4;
            173: spo = 5'h5;
            174: spo = 5'h6;
            175: spo = 5'h7;
            176: spo = 5'h19;
            177: spo = 5'h1a;
            178: spo = 5'h1b;
            179: spo = 5'h1c;
            180: spo = 5'h1d;
            181: spo = 5'h1e;
            182: spo = 5'h1f;
            183: spo = 5'h0;
            184: spo = 5'h1;
            185: spo = 5'h2;
            186: spo = 5'h2;
            187: spo = 5'h3;
            188: spo = 5'h4;
            189: spo = 5'h5;
            190: spo = 5'h6;
            191: spo = 5'h7;
            192: spo = 5'h19;
            193: spo = 5'h1a;
            194: spo = 5'h1b;
            195: spo = 5'h1c;
            196: spo = 5'h1d;
            197: spo = 5'h1e;
            198: spo = 5'h1f;
            199: spo = 5'h0;
            200: spo = 5'h1;
            201: spo = 5'h2;
            202: spo = 5'h3;
            203: spo = 5'h4;
            204: spo = 5'h5;
            205: spo = 5'h6;
            206: spo = 5'h7;
            207: spo = 5'h8;
            208: spo = 5'h19;
            209: spo = 5'h1a;
            210: spo = 5'h1b;
            211: spo = 5'h1c;
            212: spo = 5'h1d;
            213: spo = 5'h1e;
            214: spo = 5'h1f;
            215: spo = 5'h0;
            216: spo = 5'h1;
            217: spo = 5'h2;
            218: spo = 5'h3;
            219: spo = 5'h4;
            220: spo = 5'h5;
            221: spo = 5'h6;
            222: spo = 5'h7;
            223: spo = 5'h8;
            224: spo = 5'h19;
            225: spo = 5'h1a;
            226: spo = 5'h1b;
            227: spo = 5'h1c;
            228: spo = 5'h1d;
            229: spo = 5'h1e;
            230: spo = 5'h1f;
            231: spo = 5'h0;
            232: spo = 5'h1;
            233: spo = 5'h2;
            234: spo = 5'h3;
            235: spo = 5'h4;
            236: spo = 5'h5;
            237: spo = 5'h6;
            238: spo = 5'h7;
            239: spo = 5'h8;
            240: spo = 5'h19;
            241: spo = 5'h1a;
            242: spo = 5'h1b;
            243: spo = 5'h1c;
            244: spo = 5'h1d;
            245: spo = 5'h1e;
            246: spo = 5'h1f;
            247: spo = 5'h0;
            248: spo = 5'h1;
            249: spo = 5'h2;
            250: spo = 5'h3;
            251: spo = 5'h4;
            252: spo = 5'h5;
            253: spo = 5'h6;
            254: spo = 5'h7;
            255: spo = 5'h8;
            default: spo = 5'h0;
		endcase
	end
endmodule